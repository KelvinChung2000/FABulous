(* blackbox *)
module ALU #(
    parameter ALU_func = 0
)
(
    input [31:0] data_in1,
    input [31:0] data_in2,
    input [31:0] data_in3,
    output [31:0] data_out
);

endmodule
