module mults1 #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i3_data_size1;
wire[WIDTH-1:0] i3_mul1;
wire[WIDTH-1:0] i3_add1;
wire[WIDTH-1:0] i4_load;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i5_mul;
wire[WIDTH-1:0] i6_add;
wire[WIDTH-1:0] i7_data_size1;
wire[WIDTH-1:0] i7_mul1;
wire[WIDTH-1:0] i7_add1;
wire[WIDTH-1:0] i8_load;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i9_mul;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i10_add;
wire[WIDTH-1:0] i11_data_size1;
wire[WIDTH-1:0] i11_mul1;
wire[WIDTH-1:0] i11_add1;
wire[WIDTH-1:0] i12_load;
wire[WIDTH-1:0] const6;
wire[WIDTH-1:0] i13_mul;
wire[WIDTH-1:0] const7;
wire[WIDTH-1:0] i14_add;
wire[WIDTH-1:0] i15_data_size1;
wire[WIDTH-1:0] i15_mul1;
wire[WIDTH-1:0] i15_add1;
wire[WIDTH-1:0] i16_load;
wire[WIDTH-1:0] const8;
wire[WIDTH-1:0] i17_mul;
wire[WIDTH-1:0] i18_add;
wire[WIDTH-1:0] i19_add;
wire[WIDTH-1:0] i20_add;
wire[WIDTH-1:0] i21_add;
wire[WIDTH-1:0] input0;
wire i22_icmp;
wire[WIDTH-1:0] const2_dup_1;
wire[WIDTH-1:0] const2_dup_2;
wire[WIDTH-1:0] const2_dup_3;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i3_data_size1_alu;
wire[WIDTH-1:0] i3_mul1_alu;
wire[WIDTH-1:0] i3_add1_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i5_mul_alu;
wire[WIDTH-1:0] i6_add_alu;
wire[WIDTH-1:0] i7_data_size1_alu;
wire[WIDTH-1:0] i7_mul1_alu;
wire[WIDTH-1:0] i7_add1_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i9_mul_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i10_add_alu;
wire[WIDTH-1:0] i11_data_size1_alu;
wire[WIDTH-1:0] i11_mul1_alu;
wire[WIDTH-1:0] i11_add1_alu;
wire[WIDTH-1:0] const6_alu;
wire[WIDTH-1:0] i13_mul_alu;
wire[WIDTH-1:0] const7_alu;
wire[WIDTH-1:0] i14_add_alu;
wire[WIDTH-1:0] i15_data_size1_alu;
wire[WIDTH-1:0] i15_mul1_alu;
wire[WIDTH-1:0] i15_add1_alu;
wire[WIDTH-1:0] const8_alu;
wire[WIDTH-1:0] i17_mul_alu;
wire[WIDTH-1:0] i18_add_alu;
wire[WIDTH-1:0] i19_add_alu;
wire[WIDTH-1:0] i20_add_alu;
wire[WIDTH-1:0] i21_add_alu;
wire[WIDTH-1:0] i21_output_alu;
wire[WIDTH-1:0] const2_dup_1_alu;
wire[WIDTH-1:0] const2_dup_2_alu;
wire[WIDTH-1:0] const2_dup_3_alu;
wire[WIDTH-1:0] i23_br;
wire[WIDTH-1:0] i21_output;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(1)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const2(.const_out(const2));
const_unit #(.ConfigBits(4)) inst_i3_data_size1(.const_out(i3_data_size1));
ALU #(.ALU_func(mul_op)) inst_i3_mul1(.data_in1(i3_data_size1), .data_in2(i6_add), .data_in3(), .data_out(i3_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_mul1_reg(.reg_in(i3_mul1_alu), .reg_out(i3_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i3_add1(.data_in1(const2), .data_in2(i3_mul1), .data_in3(), .data_out(i3_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add1_reg(.reg_in(i3_add1_alu), .reg_out(i3_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i4_load(.addr0(i3_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i4_load));
const_unit #(.ConfigBits(10)) inst_const3(.const_out(const3));
ALU #(.ALU_func(mul_op)) inst_i5_mul(.data_in1(i4_load), .data_in2(const3), .data_in3(), .data_out(i5_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_mul_reg(.reg_in(i5_mul_alu), .reg_out(i5_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i6_add(.data_in1(const0), .data_in2(i6_add), .data_in3(), .data_out(i6_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add_reg(.reg_in(i6_add_alu), .reg_out(i6_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i7_data_size1(.const_out(i7_data_size1));
ALU #(.ALU_func(mul_op)) inst_i7_mul1(.data_in1(i6_add), .data_in2(i7_data_size1), .data_in3(), .data_out(i7_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_mul1_reg(.reg_in(i7_mul1_alu), .reg_out(i7_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i7_add1(.data_in1(i7_mul1), .data_in2(const2_dup_1), .data_in3(), .data_out(i7_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_add1_reg(.reg_in(i7_add1_alu), .reg_out(i7_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i8_load(.addr0(i7_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i8_load));
const_unit #(.ConfigBits(20)) inst_const4(.const_out(const4));
ALU #(.ALU_func(mul_op)) inst_i9_mul(.data_in1(i8_load), .data_in2(const4), .data_in3(), .data_out(i9_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_mul_reg(.reg_in(i9_mul_alu), .reg_out(i9_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2)) inst_const5(.const_out(const5));
ALU #(.ALU_func(add_op)) inst_i10_add(.data_in1(const5), .data_in2(i6_add), .data_in3(), .data_out(i10_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_add_reg(.reg_in(i10_add_alu), .reg_out(i10_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i11_data_size1(.const_out(i11_data_size1));
ALU #(.ALU_func(mul_op)) inst_i11_mul1(.data_in1(i10_add), .data_in2(i11_data_size1), .data_in3(), .data_out(i11_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_mul1_reg(.reg_in(i11_mul1_alu), .reg_out(i11_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i11_add1(.data_in1(i11_mul1), .data_in2(const2_dup_2), .data_in3(), .data_out(i11_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_add1_reg(.reg_in(i11_add1_alu), .reg_out(i11_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i12_load(.addr0(i11_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i12_load));
const_unit #(.ConfigBits(39)) inst_const6(.const_out(const6));
ALU #(.ALU_func(mul_op)) inst_i13_mul(.data_in1(i12_load), .data_in2(const6), .data_in3(), .data_out(i13_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i13_mul_reg(.reg_in(i13_mul_alu), .reg_out(i13_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(3)) inst_const7(.const_out(const7));
ALU #(.ALU_func(add_op)) inst_i14_add(.data_in1(const7), .data_in2(i6_add), .data_in3(), .data_out(i14_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_add_reg(.reg_in(i14_add_alu), .reg_out(i14_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i15_data_size1(.const_out(i15_data_size1));
ALU #(.ALU_func(mul_op)) inst_i15_mul1(.data_in1(i14_add), .data_in2(i15_data_size1), .data_in3(), .data_out(i15_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_mul1_reg(.reg_in(i15_mul1_alu), .reg_out(i15_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i15_add1(.data_in1(i15_mul1), .data_in2(const2_dup_3), .data_in3(), .data_out(i15_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_add1_reg(.reg_in(i15_add1_alu), .reg_out(i15_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i16_load(.addr0(i15_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i16_load));
const_unit #(.ConfigBits(15)) inst_const8(.const_out(const8));
ALU #(.ALU_func(mul_op)) inst_i17_mul(.data_in1(i16_load), .data_in2(const8), .data_in3(), .data_out(i17_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i17_mul_reg(.reg_in(i17_mul_alu), .reg_out(i17_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i18_add(.data_in1(i5_mul), .data_in2(i21_add), .data_in3(), .data_out(i18_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i18_add_reg(.reg_in(i18_add_alu), .reg_out(i18_add), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i19_add(.data_in1(i9_mul), .data_in2(i18_add), .data_in3(), .data_out(i19_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i19_add_reg(.reg_in(i19_add_alu), .reg_out(i19_add), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i20_add(.data_in1(i13_mul), .data_in2(i19_add), .data_in3(), .data_out(i20_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i20_add_reg(.reg_in(i20_add_alu), .reg_out(i20_add), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i21_add(.data_in1(i17_mul), .data_in2(i20_add), .data_in3(), .data_out(i21_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i21_add_reg(.reg_in(i21_add_alu), .reg_out(i21_add), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i22_icmp(.A(i6_add), .B(input0), .Y(i22_icmp));
(* keep *) IO_WIDTH_1 inst_i23_br(.from_fabric(i22_icmp), .in(), .to_fabric(), .out());
(* keep *) IO inst_i21_output(.from_fabric(i21_add), .in(), .to_fabric(), .out());
const_unit #(.ConfigBits(2560)) inst_const2_dup_1(.const_out(const2_dup_1));
const_unit #(.ConfigBits(2560)) inst_const2_dup_2(.const_out(const2_dup_2));
const_unit #(.ConfigBits(2560)) inst_const2_dup_3(.const_out(const2_dup_3));

endmodule
