module test();

  wire [31:0] in;
  wire [31:0] out;
  assign out = in + 16;

endmodule