(* blackbox *)
module IO #(
)
(
    input wire[31:0] N_from_fabric,
    input wire[31:0] N_in,
    output reg[31:0] N_to_fabric,
    output reg[31:0] N_out
);

endmodule

