module IO #() (
    (* FABulous, BUS *) input in,
    (* FABulous, BUS *) output out,
    (* FABulous, CONFIG_BIT, IO *) input ConfigBits
);
endmodule
