module matrixmultiply #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i3_data_size1;
wire[WIDTH-1:0] input0;
wire[WIDTH-1:0] i3_mul1;
wire[WIDTH-1:0] i3_add1;
wire[WIDTH-1:0] i3_mul2;
wire[WIDTH-1:0] i3_add2;
wire[WIDTH-1:0] i4_load;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i5_data_size1;
wire[WIDTH-1:0] i5_mul1;
wire[WIDTH-1:0] i5_add1;
wire[WIDTH-1:0] i5_data_size2;
wire[WIDTH-1:0] input1;
wire[WIDTH-1:0] i5_mul2;
wire[WIDTH-1:0] i5_add2;
wire[WIDTH-1:0] i6_load;
wire[WIDTH-1:0] i7_mul;
wire[WIDTH-1:0] i8_add;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i9_add;
wire[WIDTH-1:0] const5;
wire i10_icmp;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i3_data_size1_alu;
wire[WIDTH-1:0] i3_mul1_alu;
wire[WIDTH-1:0] i3_add1_alu;
wire[WIDTH-1:0] i3_mul2_alu;
wire[WIDTH-1:0] i3_add2_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i5_data_size1_alu;
wire[WIDTH-1:0] i5_mul1_alu;
wire[WIDTH-1:0] i5_add1_alu;
wire[WIDTH-1:0] i5_data_size2_alu;
wire[WIDTH-1:0] i5_mul2_alu;
wire[WIDTH-1:0] i5_add2_alu;
wire[WIDTH-1:0] i7_mul_alu;
wire[WIDTH-1:0] i8_add_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i9_add_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i8_output_alu;
wire[WIDTH-1:0] i11_br;
wire[WIDTH-1:0] i8_output;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(0)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const2(.const_out(const2));
const_unit #(.ConfigBits(80)) inst_i3_data_size1(.const_out(i3_data_size1));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
ALU #(.ALU_func(mul_op)) inst_i3_mul1(.data_in1(i3_data_size1), .data_in2(input0), .data_in3(), .data_out(i3_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_mul1_reg(.reg_in(i3_mul1_alu), .reg_out(i3_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i3_add1(.data_in1(const2), .data_in2(i3_mul1), .data_in3(), .data_out(i3_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add1_reg(.reg_in(i3_add1_alu), .reg_out(i3_add1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i3_mul2(.data_in1(const0), .data_in2(i9_add), .data_in3(), .data_out(i3_mul2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_mul2_reg(.reg_in(i3_mul2_alu), .reg_out(i3_mul2), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i3_add2(.data_in1(i3_add1), .data_in2(i3_mul2), .data_in3(), .data_out(i3_add2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add2_reg(.reg_in(i3_add2_alu), .reg_out(i3_add2), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i4_load(.addr0(i3_add2), .reset(global_rst), .write_data(), .write_en(), .read_data(i4_load));
const_unit #(.ConfigBits(2816)) inst_const3(.const_out(const3));
const_unit #(.ConfigBits(80)) inst_i5_data_size1(.const_out(i5_data_size1));
ALU #(.ALU_func(mul_op)) inst_i5_mul1(.data_in1(i5_data_size1), .data_in2(i9_add), .data_in3(), .data_out(i5_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_mul1_reg(.reg_in(i5_mul1_alu), .reg_out(i5_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i5_add1(.data_in1(const3), .data_in2(i5_mul1), .data_in3(), .data_out(i5_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_add1_reg(.reg_in(i5_add1_alu), .reg_out(i5_add1), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i5_data_size2(.const_out(i5_data_size2));
(* keep *) IO inst_input1(.from_fabric(), .in(), .to_fabric(input1), .out());
ALU #(.ALU_func(mul_op)) inst_i5_mul2(.data_in1(i5_data_size2), .data_in2(input1), .data_in3(), .data_out(i5_mul2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_mul2_reg(.reg_in(i5_mul2_alu), .reg_out(i5_mul2), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i5_add2(.data_in1(i5_add1), .data_in2(i5_mul2), .data_in3(), .data_out(i5_add2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_add2_reg(.reg_in(i5_add2_alu), .reg_out(i5_add2), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i6_load(.addr0(i5_add2), .reset(global_rst), .write_data(), .write_en(), .read_data(i6_load));
ALU #(.ALU_func(mul_op)) inst_i7_mul(.data_in1(i4_load), .data_in2(i6_load), .data_in3(), .data_out(i7_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_mul_reg(.reg_in(i7_mul_alu), .reg_out(i7_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i8_add(.data_in1(i7_mul), .data_in2(i8_add), .data_in3(), .data_out(i8_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_add_reg(.reg_in(i8_add_alu), .reg_out(i8_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(1)) inst_const4(.const_out(const4));
ALU #(.ALU_func(add_op)) inst_i9_add(.data_in1(const4), .data_in2(i9_add), .data_in3(), .data_out(i9_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add_reg(.reg_in(i9_add_alu), .reg_out(i9_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(20)) inst_const5(.const_out(const5));
compare #(.conf(0)) inst_i10_icmp(.A(i9_add), .B(const5), .Y(i10_icmp));
(* keep *) IO_WIDTH_1 inst_i11_br(.from_fabric(i10_icmp), .in(), .to_fabric(), .out());
(* keep *) IO inst_i8_output(.from_fabric(i8_add), .in(), .to_fabric(), .out());

endmodule
