module handshake_buffer_2slots_seq_1ins_1outs_ctrl (
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0_valid
);
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			ready0_reg <= 1'h0;
			valid1_reg <= 1'h0;
			ready1_reg <= 1'h0;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			ready0_reg <= ~(_GEN_0 & ready0_reg) & (~_GEN_0 & ~ready0_reg ? valid0_reg : ready0_reg);
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			ready1_reg <= ~(out0_ready & ready1_reg) & (~out0_ready & ~ready1_reg ? valid1_reg : ready1_reg);
		end
	assign in0_ready = _GEN;
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module handshake_buffer_in_ui32_out_ui32_2slots_seq (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input [31:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg [31:0] data0_reg;
	reg [31:0] ctrl_data0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	reg [31:0] data1_reg;
	reg [31:0] ctrl_data1_reg;
	wire _GEN_1 = ~_GEN_0 & ~ready0_reg;
	wire _GEN_2 = _GEN_0 & ready0_reg;
	wire _GEN_3 = ~out0_ready & ~ready1_reg;
	wire _GEN_4 = out0_ready & ready1_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			data0_reg <= 32'h00000000;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= 32'h00000000;
			valid1_reg <= 1'h0;
			data1_reg <= 32'h00000000;
			ready1_reg <= 1'h0;
			ctrl_data1_reg <= 32'h00000000;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_2 & (_GEN_1 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= (_GEN_2 ? 32'h00000000 : (_GEN_1 ? data0_reg : ctrl_data0_reg));
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			data1_reg <= (_GEN_0 ? (ready0_reg ? ctrl_data0_reg : data0_reg) : data1_reg);
			ready1_reg <= ~_GEN_4 & (_GEN_3 ? valid1_reg : ready1_reg);
			ctrl_data1_reg <= (_GEN_4 ? 32'h00000000 : (_GEN_3 ? data1_reg : ctrl_data1_reg));
		end
	assign in0_ready = _GEN;
	assign out0 = (ready1_reg ? ctrl_data1_reg : data1_reg);
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module handshake_fork_1ins_4outs_ctrl (
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	in0_ready,
	out0_valid,
	out1_valid,
	out2_valid,
	out3_valid
);
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	output wire in0_ready;
	output wire out0_valid;
	output wire out1_valid;
	output wire out2_valid;
	output wire out3_valid;
	wire allDone;
	wire done3;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
		end
	wire _GEN_2 = ~emitted_3 & in0_valid;
	assign done3 = (out3_ready & _GEN_2) | emitted_3;
	assign allDone = ((done0 & done1) & done2) & done3;
	assign in0_ready = allDone;
	assign out0_valid = _GEN;
	assign out1_valid = _GEN_0;
	assign out2_valid = _GEN_1;
	assign out3_valid = _GEN_2;
endmodule
module handshake_fork_in_ui32_out_ui32_ui32 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid
);
	input [31:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	output wire in0_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	output wire [31:0] out1;
	output wire out1_valid;
	wire allDone;
	wire done1;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
		end
	wire _GEN_0 = ~emitted_1 & in0_valid;
	assign done1 = (out1_ready & _GEN_0) | emitted_1;
	assign allDone = done0 & done1;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
endmodule
module handshake_join_in_ui32_1ins_1outs_ctrl (
	in0,
	in0_valid,
	out0_ready,
	in0_ready,
	out0_valid
);
	input [31:0] in0;
	input in0_valid;
	input out0_ready;
	output wire in0_ready;
	output wire out0_valid;
	assign in0_ready = out0_ready & in0_valid;
	assign out0_valid = in0_valid;
endmodule
module arith_index_cast_in_ui64_out_ui10 (
	in0,
	in0_valid,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input [63:0] in0;
	input in0_valid;
	input out0_ready;
	output wire in0_ready;
	output wire [9:0] out0;
	output wire out0_valid;
	assign in0_ready = out0_ready & in0_valid;
	assign out0 = in0[9:0];
	assign out0_valid = in0_valid;
endmodule
module handshake_buffer_in_ui10_out_ui10_2slots_seq (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input [9:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire [9:0] out0;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg [9:0] data0_reg;
	reg [9:0] ctrl_data0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	reg [9:0] data1_reg;
	reg [9:0] ctrl_data1_reg;
	wire _GEN_1 = ~_GEN_0 & ~ready0_reg;
	wire _GEN_2 = _GEN_0 & ready0_reg;
	wire _GEN_3 = ~out0_ready & ~ready1_reg;
	wire _GEN_4 = out0_ready & ready1_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			data0_reg <= 10'h000;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= 10'h000;
			valid1_reg <= 1'h0;
			data1_reg <= 10'h000;
			ready1_reg <= 1'h0;
			ctrl_data1_reg <= 10'h000;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_2 & (_GEN_1 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= (_GEN_2 ? 10'h000 : (_GEN_1 ? data0_reg : ctrl_data0_reg));
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			data1_reg <= (_GEN_0 ? (ready0_reg ? ctrl_data0_reg : data0_reg) : data1_reg);
			ready1_reg <= ~_GEN_4 & (_GEN_3 ? valid1_reg : ready1_reg);
			ctrl_data1_reg <= (_GEN_4 ? 10'h000 : (_GEN_3 ? data1_reg : ctrl_data1_reg));
		end
	assign in0_ready = _GEN;
	assign out0 = (ready1_reg ? ctrl_data1_reg : data1_reg);
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module hw_struct_create_in_ui10_ui32_out_struct_address_ui10_data_ui32 (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [9:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [41:0] out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = {in0, in1};
	assign out0_valid = _GEN;
endmodule
module handshake_buffer_in_struct_address_ui10_data_ui32_out_struct_address_ui10_data_ui32_2slots_seq (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input wire [41:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire [41:0] out0;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg [41:0] data0_reg;
	reg [41:0] ctrl_data0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	reg [41:0] data1_reg;
	reg [41:0] ctrl_data1_reg;
	wire [41:0] _GEN_1 = 42'h00000000000;
	wire _GEN_2 = ~_GEN_0 & ~ready0_reg;
	wire _GEN_3 = _GEN_0 & ready0_reg;
	wire _GEN_4 = ~out0_ready & ~ready1_reg;
	wire _GEN_5 = out0_ready & ready1_reg;
	wire [41:0] _GEN_6 = 42'h00000000000;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			data0_reg <= _GEN_6;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= _GEN_6;
			valid1_reg <= 1'h0;
			data1_reg <= _GEN_6;
			ready1_reg <= 1'h0;
			ctrl_data1_reg <= _GEN_6;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_3 & (_GEN_2 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= (_GEN_3 ? _GEN_1 : (_GEN_2 ? data0_reg : ctrl_data0_reg));
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			data1_reg <= (_GEN_0 ? (ready0_reg ? ctrl_data0_reg : data0_reg) : data1_reg);
			ready1_reg <= ~_GEN_5 & (_GEN_4 ? valid1_reg : ready1_reg);
			ctrl_data1_reg <= (_GEN_5 ? _GEN_1 : (_GEN_4 ? data1_reg : ctrl_data1_reg));
		end
	assign in0_ready = _GEN;
	assign out0 = (ready1_reg ? ctrl_data1_reg : data1_reg);
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module handshake_constant_c0_out_ui64 (
	ctrl_valid,
	out0_ready,
	ctrl_ready,
	out0,
	out0_valid
);
	input ctrl_valid;
	input out0_ready;
	output wire ctrl_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	assign ctrl_ready = out0_ready;
	assign out0 = 64'h0000000000000000;
	assign out0_valid = ctrl_valid;
endmodule
module handshake_buffer_in_ui64_out_ui64_2slots_seq (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input [63:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg [63:0] data0_reg;
	reg [63:0] ctrl_data0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	reg [63:0] data1_reg;
	reg [63:0] ctrl_data1_reg;
	wire _GEN_1 = ~_GEN_0 & ~ready0_reg;
	wire _GEN_2 = _GEN_0 & ready0_reg;
	wire _GEN_3 = ~out0_ready & ~ready1_reg;
	wire _GEN_4 = out0_ready & ready1_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			data0_reg <= 64'h0000000000000000;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= 64'h0000000000000000;
			valid1_reg <= 1'h0;
			data1_reg <= 64'h0000000000000000;
			ready1_reg <= 1'h0;
			ctrl_data1_reg <= 64'h0000000000000000;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_2 & (_GEN_1 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= (_GEN_2 ? 64'h0000000000000000 : (_GEN_1 ? data0_reg : ctrl_data0_reg));
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			data1_reg <= (_GEN_0 ? (ready0_reg ? ctrl_data0_reg : data0_reg) : data1_reg);
			ready1_reg <= ~_GEN_4 & (_GEN_3 ? valid1_reg : ready1_reg);
			ctrl_data1_reg <= (_GEN_4 ? 64'h0000000000000000 : (_GEN_3 ? data1_reg : ctrl_data1_reg));
		end
	assign in0_ready = _GEN;
	assign out0 = (ready1_reg ? ctrl_data1_reg : data1_reg);
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module handshake_constant_c20_out_ui64 (
	ctrl_valid,
	out0_ready,
	ctrl_ready,
	out0,
	out0_valid
);
	input ctrl_valid;
	input out0_ready;
	output wire ctrl_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	assign ctrl_ready = out0_ready;
	assign out0 = 64'h0000000000000014;
	assign out0_valid = ctrl_valid;
endmodule
module handshake_constant_c1_out_ui64 (
	ctrl_valid,
	out0_ready,
	ctrl_ready,
	out0,
	out0_valid
);
	input ctrl_valid;
	input out0_ready;
	output wire ctrl_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	assign ctrl_ready = out0_ready;
	assign out0 = 64'h0000000000000001;
	assign out0_valid = ctrl_valid;
endmodule
module handshake_buffer_in_ui1_out_ui1_1slots_seq_init_0 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg data0_reg;
	reg ctrl_data0_reg;
	wire _GEN_0 = ~out0_ready & ~ready0_reg;
	wire _GEN_1 = out0_ready & ready0_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h1;
			data0_reg <= 1'h0;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= 1'h0;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_1 & (_GEN_0 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= ~_GEN_1 & (_GEN_0 ? data0_reg : ctrl_data0_reg);
		end
	assign in0_ready = _GEN;
	assign out0 = (ready0_reg ? ctrl_data0_reg : data0_reg);
	assign out0_valid = (ready0_reg ? ready0_reg : valid0_reg);
endmodule
module handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	output wire out1;
	output wire out1_valid;
	output wire out2;
	output wire out2_valid;
	output wire out3;
	output wire out3_valid;
	output wire out4;
	output wire out4_valid;
	output wire out5;
	output wire out5_valid;
	wire allDone;
	wire done5;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
		end
	wire _GEN_4 = ~emitted_5 & in0_valid;
	assign done5 = (out5_ready & _GEN_4) | emitted_5;
	assign allDone = ((((done0 & done1) & done2) & done3) & done4) & done5;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
endmodule
module handshake_buffer_in_ui1_out_ui1_2slots_seq (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	in0_ready,
	out0,
	out0_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	reg ready1_reg;
	reg ready0_reg;
	reg valid0_reg;
	wire _GEN = ~valid0_reg | ~ready0_reg;
	reg data0_reg;
	reg ctrl_data0_reg;
	reg valid1_reg;
	wire _GEN_0 = ~valid1_reg | ~ready1_reg;
	reg data1_reg;
	reg ctrl_data1_reg;
	wire _GEN_1 = ~_GEN_0 & ~ready0_reg;
	wire _GEN_2 = _GEN_0 & ready0_reg;
	wire _GEN_3 = ~out0_ready & ~ready1_reg;
	wire _GEN_4 = out0_ready & ready1_reg;
	always @(posedge clock)
		if (reset) begin
			valid0_reg <= 1'h0;
			data0_reg <= 1'h0;
			ready0_reg <= 1'h0;
			ctrl_data0_reg <= 1'h0;
			valid1_reg <= 1'h0;
			data1_reg <= 1'h0;
			ready1_reg <= 1'h0;
			ctrl_data1_reg <= 1'h0;
		end
		else begin
			valid0_reg <= (_GEN ? in0_valid : valid0_reg);
			data0_reg <= (_GEN ? in0 : data0_reg);
			ready0_reg <= ~_GEN_2 & (_GEN_1 ? valid0_reg : ready0_reg);
			ctrl_data0_reg <= ~_GEN_2 & (_GEN_1 ? data0_reg : ctrl_data0_reg);
			valid1_reg <= (_GEN_0 ? (ready0_reg ? ready0_reg : valid0_reg) : valid1_reg);
			data1_reg <= (_GEN_0 ? (ready0_reg ? ctrl_data0_reg : data0_reg) : data1_reg);
			ready1_reg <= ~_GEN_4 & (_GEN_3 ? valid1_reg : ready1_reg);
			ctrl_data1_reg <= ~_GEN_4 & (_GEN_3 ? data1_reg : ctrl_data1_reg);
		end
	assign in0_ready = _GEN;
	assign out0 = (ready1_reg ? ctrl_data1_reg : data1_reg);
	assign out0_valid = (ready1_reg ? ready1_reg : valid1_reg);
endmodule
module handshake_mux_in_ui1_3ins_1outs_ctrl (
	select,
	select_valid,
	in0_valid,
	in1_valid,
	out0_ready,
	select_ready,
	in0_ready,
	in1_ready,
	out0_valid
);
	input select;
	input select_valid;
	input in0_valid;
	input in1_valid;
	input out0_ready;
	output wire select_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire out0_valid;
	wire [1:0] _GEN = 2'h1 << select;
	wire _GEN_0 = (select ? in1_valid : in0_valid) & select_valid;
	wire _GEN_1 = _GEN_0 & out0_ready;
	assign select_ready = _GEN_1;
	assign in0_ready = _GEN[0] & _GEN_1;
	assign in1_ready = _GEN[1] & _GEN_1;
	assign out0_valid = _GEN_0;
endmodule
module handshake_mux_in_ui1_ui64_ui64_out_ui64 (
	select,
	select_valid,
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	select_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input select;
	input select_valid;
	input [63:0] in0;
	input in0_valid;
	input [63:0] in1;
	input in1_valid;
	input out0_ready;
	output wire select_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	wire [1:0] _GEN = 2'h1 << select;
	wire _GEN_0 = (select ? in1_valid : in0_valid) & select_valid;
	wire _GEN_1 = _GEN_0 & out0_ready;
	assign select_ready = _GEN_1;
	assign in0_ready = _GEN[0] & _GEN_1;
	assign in1_ready = _GEN[1] & _GEN_1;
	assign out0 = (select ? in1 : in0);
	assign out0_valid = _GEN_0;
endmodule
module handshake_fork_in_ui64_out_ui64_ui64 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid
);
	input [63:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	output wire in0_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	output wire [63:0] out1;
	output wire out1_valid;
	wire allDone;
	wire done1;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
		end
	wire _GEN_0 = ~emitted_1 & in0_valid;
	assign done1 = (out1_ready & _GEN_0) | emitted_1;
	assign allDone = done0 & done1;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
endmodule
module handshake_mux_in_ui1_ui32_ui32_out_ui32 (
	select,
	select_valid,
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	select_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input select;
	input select_valid;
	input [31:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input out0_ready;
	output wire select_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	wire [1:0] _GEN = 2'h1 << select;
	wire _GEN_0 = (select ? in1_valid : in0_valid) & select_valid;
	wire _GEN_1 = _GEN_0 & out0_ready;
	assign select_ready = _GEN_1;
	assign in0_ready = _GEN[0] & _GEN_1;
	assign in1_ready = _GEN[1] & _GEN_1;
	assign out0 = (select ? in1 : in0);
	assign out0_valid = _GEN_0;
endmodule
module arith_cmpi_in_ui64_ui64_out_ui1_slt (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [63:0] in0;
	input in0_valid;
	input [63:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = $signed(in0) < $signed(in1);
	assign out0_valid = _GEN;
endmodule
module handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	out6_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid,
	out6,
	out6_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	input out6_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	output wire out1;
	output wire out1_valid;
	output wire out2;
	output wire out2_valid;
	output wire out3;
	output wire out3_valid;
	output wire out4;
	output wire out4_valid;
	output wire out5;
	output wire out5_valid;
	output wire out6;
	output wire out6_valid;
	wire allDone;
	wire done6;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	wire _GEN_4 = ~emitted_5 & in0_valid;
	wire done5 = (out5_ready & _GEN_4) | emitted_5;
	reg emitted_6;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
			emitted_6 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
			emitted_6 <= done6 & ~allDone;
		end
	wire _GEN_5 = ~emitted_6 & in0_valid;
	assign done6 = (out6_ready & _GEN_5) | emitted_6;
	assign allDone = (((((done0 & done1) & done2) & done3) & done4) & done5) & done6;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
	assign out6 = in0;
	assign out6_valid = _GEN_5;
endmodule
module handshake_cond_br_in_ui1_ui64_out_ui64_ui64 (
	cond,
	cond_valid,
	data,
	data_valid,
	outTrue_ready,
	outFalse_ready,
	cond_ready,
	data_ready,
	outTrue,
	outTrue_valid,
	outFalse,
	outFalse_valid
);
	input cond;
	input cond_valid;
	input [63:0] data;
	input data_valid;
	input outTrue_ready;
	input outFalse_ready;
	output wire cond_ready;
	output wire data_ready;
	output wire [63:0] outTrue;
	output wire outTrue_valid;
	output wire [63:0] outFalse;
	output wire outFalse_valid;
	wire _GEN = cond_valid & data_valid;
	wire _GEN_0 = (cond ? outTrue_ready : outFalse_ready) & _GEN;
	assign cond_ready = _GEN_0;
	assign data_ready = _GEN_0;
	assign outTrue = data;
	assign outTrue_valid = cond & _GEN;
	assign outFalse = data;
	assign outFalse_valid = ~cond & _GEN;
endmodule
module handshake_sink_in_ui64 (
	in0,
	in0_valid,
	in0_ready
);
	input [63:0] in0;
	input in0_valid;
	output wire in0_ready;
	assign in0_ready = 1'h1;
endmodule
module handshake_cond_br_in_ui1_ui32_out_ui32_ui32 (
	cond,
	cond_valid,
	data,
	data_valid,
	outTrue_ready,
	outFalse_ready,
	cond_ready,
	data_ready,
	outTrue,
	outTrue_valid,
	outFalse,
	outFalse_valid
);
	input cond;
	input cond_valid;
	input [31:0] data;
	input data_valid;
	input outTrue_ready;
	input outFalse_ready;
	output wire cond_ready;
	output wire data_ready;
	output wire [31:0] outTrue;
	output wire outTrue_valid;
	output wire [31:0] outFalse;
	output wire outFalse_valid;
	wire _GEN = cond_valid & data_valid;
	wire _GEN_0 = (cond ? outTrue_ready : outFalse_ready) & _GEN;
	assign cond_ready = _GEN_0;
	assign data_ready = _GEN_0;
	assign outTrue = data;
	assign outTrue_valid = cond & _GEN;
	assign outFalse = data;
	assign outFalse_valid = ~cond & _GEN;
endmodule
module handshake_sink_in_ui32 (
	in0,
	in0_valid,
	in0_ready
);
	input [31:0] in0;
	input in0_valid;
	output wire in0_ready;
	assign in0_ready = 1'h1;
endmodule
module handshake_cond_br_in_ui1_2ins_2outs_ctrl (
	cond,
	cond_valid,
	data_valid,
	outTrue_ready,
	outFalse_ready,
	cond_ready,
	data_ready,
	outTrue_valid,
	outFalse_valid
);
	input cond;
	input cond_valid;
	input data_valid;
	input outTrue_ready;
	input outFalse_ready;
	output wire cond_ready;
	output wire data_ready;
	output wire outTrue_valid;
	output wire outFalse_valid;
	wire _GEN = cond_valid & data_valid;
	wire _GEN_0 = (cond ? outTrue_ready : outFalse_ready) & _GEN;
	assign cond_ready = _GEN_0;
	assign data_ready = _GEN_0;
	assign outTrue_valid = cond & _GEN;
	assign outFalse_valid = ~cond & _GEN;
endmodule
module handshake_mux_in_ui64_ui64_ui64_out_ui64 (
	select,
	select_valid,
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	select_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [63:0] select;
	input select_valid;
	input [63:0] in0;
	input in0_valid;
	input [63:0] in1;
	input in1_valid;
	input out0_ready;
	output wire select_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	wire [1:0] _GEN = 2'h1 << select[0];
	wire _GEN_0 = (select[0] ? in1_valid : in0_valid) & select_valid;
	wire _GEN_1 = _GEN_0 & out0_ready;
	assign select_ready = _GEN_1;
	assign in0_ready = _GEN[0] & _GEN_1;
	assign in1_ready = _GEN[1] & _GEN_1;
	assign out0 = (select[0] ? in1 : in0);
	assign out0_valid = _GEN_0;
endmodule
module handshake_mux_in_ui64_ui32_ui32_out_ui32 (
	select,
	select_valid,
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	select_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [63:0] select;
	input select_valid;
	input [31:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input out0_ready;
	output wire select_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	wire [1:0] _GEN = 2'h1 << select[0];
	wire _GEN_0 = (select[0] ? in1_valid : in0_valid) & select_valid;
	wire _GEN_1 = _GEN_0 & out0_ready;
	assign select_ready = _GEN_1;
	assign in0_ready = _GEN[0] & _GEN_1;
	assign in1_ready = _GEN[1] & _GEN_1;
	assign out0 = (select[0] ? in1 : in0);
	assign out0_valid = _GEN_0;
endmodule
module handshake_control_merge_out_ui64_2ins_2outs_ctrl (
	in0_valid,
	in1_valid,
	clock,
	reset,
	dataOut_ready,
	index_ready,
	in0_ready,
	in1_ready,
	dataOut_valid,
	index,
	index_valid
);
	input in0_valid;
	input in1_valid;
	input clock;
	input reset;
	input dataOut_ready;
	input index_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire dataOut_valid;
	output wire [63:0] index;
	output wire index_valid;
	wire _GEN;
	wire _GEN_0;
	wire _GEN_1;
	wire [1:0] _GEN_2;
	reg [1:0] won_reg;
	reg result_emitted_reg;
	reg index_emitted_reg;
	always @(posedge clock)
		if (reset) begin
			won_reg <= 2'h0;
			result_emitted_reg <= 1'h0;
			index_emitted_reg <= 1'h0;
		end
		else begin
			won_reg <= (_GEN ? 2'h0 : _GEN_2);
			result_emitted_reg <= ~_GEN & _GEN_1;
			index_emitted_reg <= ~_GEN & _GEN_0;
		end
	assign _GEN_2 = (|won_reg ? won_reg : (in0_valid ? 2'h1 : {in1_valid, 1'h0}));
	wire _GEN_3 = |_GEN_2 & ~result_emitted_reg;
	wire _GEN_4 = |_GEN_2 & ~index_emitted_reg;
	assign _GEN_1 = (_GEN_3 & dataOut_ready) | result_emitted_reg;
	assign _GEN_0 = (_GEN_4 & index_ready) | index_emitted_reg;
	assign _GEN = _GEN_1 & _GEN_0;
	wire [1:0] _GEN_5 = (_GEN ? _GEN_2 : 2'h0);
	assign in0_ready = _GEN_5 == 2'h1;
	assign in1_ready = _GEN_5 == 2'h2;
	assign dataOut_valid = _GEN_3;
	assign index = {63'h0000000000000000, _GEN_2[1]};
	assign index_valid = _GEN_4;
endmodule
module handshake_fork_in_ui64_out_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	out6_ready,
	out7_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid,
	out6,
	out6_valid,
	out7,
	out7_valid
);
	input [63:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	input out6_ready;
	input out7_ready;
	output wire in0_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	output wire [63:0] out1;
	output wire out1_valid;
	output wire [63:0] out2;
	output wire out2_valid;
	output wire [63:0] out3;
	output wire out3_valid;
	output wire [63:0] out4;
	output wire out4_valid;
	output wire [63:0] out5;
	output wire out5_valid;
	output wire [63:0] out6;
	output wire out6_valid;
	output wire [63:0] out7;
	output wire out7_valid;
	wire allDone;
	wire done7;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	wire _GEN_4 = ~emitted_5 & in0_valid;
	wire done5 = (out5_ready & _GEN_4) | emitted_5;
	reg emitted_6;
	wire _GEN_5 = ~emitted_6 & in0_valid;
	wire done6 = (out6_ready & _GEN_5) | emitted_6;
	reg emitted_7;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
			emitted_6 <= 1'h0;
			emitted_7 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
			emitted_6 <= done6 & ~allDone;
			emitted_7 <= done7 & ~allDone;
		end
	wire _GEN_6 = ~emitted_7 & in0_valid;
	assign done7 = (out7_ready & _GEN_6) | emitted_7;
	assign allDone = ((((((done0 & done1) & done2) & done3) & done4) & done5) & done6) & done7;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
	assign out6 = in0;
	assign out6_valid = _GEN_5;
	assign out7 = in0;
	assign out7_valid = _GEN_6;
endmodule
module handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	out6_ready,
	out7_ready,
	out8_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid,
	out6,
	out6_valid,
	out7,
	out7_valid,
	out8,
	out8_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	input out6_ready;
	input out7_ready;
	input out8_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	output wire out1;
	output wire out1_valid;
	output wire out2;
	output wire out2_valid;
	output wire out3;
	output wire out3_valid;
	output wire out4;
	output wire out4_valid;
	output wire out5;
	output wire out5_valid;
	output wire out6;
	output wire out6_valid;
	output wire out7;
	output wire out7_valid;
	output wire out8;
	output wire out8_valid;
	wire allDone;
	wire done8;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	wire _GEN_4 = ~emitted_5 & in0_valid;
	wire done5 = (out5_ready & _GEN_4) | emitted_5;
	reg emitted_6;
	wire _GEN_5 = ~emitted_6 & in0_valid;
	wire done6 = (out6_ready & _GEN_5) | emitted_6;
	reg emitted_7;
	wire _GEN_6 = ~emitted_7 & in0_valid;
	wire done7 = (out7_ready & _GEN_6) | emitted_7;
	reg emitted_8;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
			emitted_6 <= 1'h0;
			emitted_7 <= 1'h0;
			emitted_8 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
			emitted_6 <= done6 & ~allDone;
			emitted_7 <= done7 & ~allDone;
			emitted_8 <= done8 & ~allDone;
		end
	wire _GEN_7 = ~emitted_8 & in0_valid;
	assign done8 = (out8_ready & _GEN_7) | emitted_8;
	assign allDone = (((((((done0 & done1) & done2) & done3) & done4) & done5) & done6) & done7) & done8;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
	assign out6 = in0;
	assign out6_valid = _GEN_5;
	assign out7 = in0;
	assign out7_valid = _GEN_6;
	assign out8 = in0;
	assign out8_valid = _GEN_7;
endmodule
module handshake_fork_1ins_6outs_ctrl (
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	in0_ready,
	out0_valid,
	out1_valid,
	out2_valid,
	out3_valid,
	out4_valid,
	out5_valid
);
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	output wire in0_ready;
	output wire out0_valid;
	output wire out1_valid;
	output wire out2_valid;
	output wire out3_valid;
	output wire out4_valid;
	output wire out5_valid;
	wire allDone;
	wire done5;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
		end
	wire _GEN_4 = ~emitted_5 & in0_valid;
	assign done5 = (out5_ready & _GEN_4) | emitted_5;
	assign allDone = ((((done0 & done1) & done2) & done3) & done4) & done5;
	assign in0_ready = allDone;
	assign out0_valid = _GEN;
	assign out1_valid = _GEN_0;
	assign out2_valid = _GEN_1;
	assign out3_valid = _GEN_2;
	assign out4_valid = _GEN_3;
	assign out5_valid = _GEN_4;
endmodule
module handshake_join_2ins_1outs_ctrl (
	in0_valid,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0_valid
);
	input in0_valid;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0_valid = _GEN;
endmodule
module handshake_constant_c30_out_ui64 (
	ctrl_valid,
	out0_ready,
	ctrl_ready,
	out0,
	out0_valid
);
	input ctrl_valid;
	input out0_ready;
	output wire ctrl_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	assign ctrl_ready = out0_ready;
	assign out0 = 64'h000000000000001e;
	assign out0_valid = ctrl_valid;
endmodule
module arith_muli_in_ui64_ui64_out_ui64 (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [63:0] in0;
	input in0_valid;
	input [63:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = in0 * in1;
	assign out0_valid = _GEN;
endmodule
module arith_addi_in_ui64_ui64_out_ui64 (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [63:0] in0;
	input in0_valid;
	input [63:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = in0 + in1;
	assign out0_valid = _GEN;
endmodule
module handshake_load_in_ui64_ui32_out_ui32_ui64 (
	addrIn0,
	addrIn0_valid,
	dataFromMem,
	dataFromMem_valid,
	ctrl_valid,
	dataOut_ready,
	addrOut0_ready,
	addrIn0_ready,
	dataFromMem_ready,
	ctrl_ready,
	dataOut,
	dataOut_valid,
	addrOut0,
	addrOut0_valid
);
	input [63:0] addrIn0;
	input addrIn0_valid;
	input [31:0] dataFromMem;
	input dataFromMem_valid;
	input ctrl_valid;
	input dataOut_ready;
	input addrOut0_ready;
	output wire addrIn0_ready;
	output wire dataFromMem_ready;
	output wire ctrl_ready;
	output wire [31:0] dataOut;
	output wire dataOut_valid;
	output wire [63:0] addrOut0;
	output wire addrOut0_valid;
	wire _GEN = addrIn0_valid & ctrl_valid;
	wire _GEN_0 = addrOut0_ready & _GEN;
	assign addrIn0_ready = _GEN_0;
	assign dataFromMem_ready = dataOut_ready;
	assign ctrl_ready = _GEN_0;
	assign dataOut = dataFromMem;
	assign dataOut_valid = dataFromMem_valid;
	assign addrOut0 = addrIn0;
	assign addrOut0_valid = _GEN;
endmodule
module arith_muli_in_ui32_ui32_out_ui32 (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [31:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = in0 * in1;
	assign out0_valid = _GEN;
endmodule
module handshake_fork_in_ui64_out_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	out6_ready,
	out7_ready,
	out8_ready,
	out9_ready,
	out10_ready,
	out11_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid,
	out6,
	out6_valid,
	out7,
	out7_valid,
	out8,
	out8_valid,
	out9,
	out9_valid,
	out10,
	out10_valid,
	out11,
	out11_valid
);
	input [63:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	input out6_ready;
	input out7_ready;
	input out8_ready;
	input out9_ready;
	input out10_ready;
	input out11_ready;
	output wire in0_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	output wire [63:0] out1;
	output wire out1_valid;
	output wire [63:0] out2;
	output wire out2_valid;
	output wire [63:0] out3;
	output wire out3_valid;
	output wire [63:0] out4;
	output wire out4_valid;
	output wire [63:0] out5;
	output wire out5_valid;
	output wire [63:0] out6;
	output wire out6_valid;
	output wire [63:0] out7;
	output wire out7_valid;
	output wire [63:0] out8;
	output wire out8_valid;
	output wire [63:0] out9;
	output wire out9_valid;
	output wire [63:0] out10;
	output wire out10_valid;
	output wire [63:0] out11;
	output wire out11_valid;
	wire allDone;
	wire done11;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	wire _GEN_4 = ~emitted_5 & in0_valid;
	wire done5 = (out5_ready & _GEN_4) | emitted_5;
	reg emitted_6;
	wire _GEN_5 = ~emitted_6 & in0_valid;
	wire done6 = (out6_ready & _GEN_5) | emitted_6;
	reg emitted_7;
	wire _GEN_6 = ~emitted_7 & in0_valid;
	wire done7 = (out7_ready & _GEN_6) | emitted_7;
	reg emitted_8;
	wire _GEN_7 = ~emitted_8 & in0_valid;
	wire done8 = (out8_ready & _GEN_7) | emitted_8;
	reg emitted_9;
	wire _GEN_8 = ~emitted_9 & in0_valid;
	wire done9 = (out9_ready & _GEN_8) | emitted_9;
	reg emitted_10;
	wire _GEN_9 = ~emitted_10 & in0_valid;
	wire done10 = (out10_ready & _GEN_9) | emitted_10;
	reg emitted_11;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
			emitted_6 <= 1'h0;
			emitted_7 <= 1'h0;
			emitted_8 <= 1'h0;
			emitted_9 <= 1'h0;
			emitted_10 <= 1'h0;
			emitted_11 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
			emitted_6 <= done6 & ~allDone;
			emitted_7 <= done7 & ~allDone;
			emitted_8 <= done8 & ~allDone;
			emitted_9 <= done9 & ~allDone;
			emitted_10 <= done10 & ~allDone;
			emitted_11 <= done11 & ~allDone;
		end
	wire _GEN_10 = ~emitted_11 & in0_valid;
	assign done11 = (out11_ready & _GEN_10) | emitted_11;
	assign allDone = ((((((((((done0 & done1) & done2) & done3) & done4) & done5) & done6) & done7) & done8) & done9) & done10) & done11;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
	assign out6 = in0;
	assign out6_valid = _GEN_5;
	assign out7 = in0;
	assign out7_valid = _GEN_6;
	assign out8 = in0;
	assign out8_valid = _GEN_7;
	assign out9 = in0;
	assign out9_valid = _GEN_8;
	assign out10 = in0;
	assign out10_valid = _GEN_9;
	assign out11 = in0;
	assign out11_valid = _GEN_10;
endmodule
module handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	out5_ready,
	out6_ready,
	out7_ready,
	out8_ready,
	out9_ready,
	out10_ready,
	out11_ready,
	out12_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid,
	out3,
	out3_valid,
	out4,
	out4_valid,
	out5,
	out5_valid,
	out6,
	out6_valid,
	out7,
	out7_valid,
	out8,
	out8_valid,
	out9,
	out9_valid,
	out10,
	out10_valid,
	out11,
	out11_valid,
	out12,
	out12_valid
);
	input in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	input out5_ready;
	input out6_ready;
	input out7_ready;
	input out8_ready;
	input out9_ready;
	input out10_ready;
	input out11_ready;
	input out12_ready;
	output wire in0_ready;
	output wire out0;
	output wire out0_valid;
	output wire out1;
	output wire out1_valid;
	output wire out2;
	output wire out2_valid;
	output wire out3;
	output wire out3_valid;
	output wire out4;
	output wire out4_valid;
	output wire out5;
	output wire out5_valid;
	output wire out6;
	output wire out6_valid;
	output wire out7;
	output wire out7_valid;
	output wire out8;
	output wire out8_valid;
	output wire out9;
	output wire out9_valid;
	output wire out10;
	output wire out10_valid;
	output wire out11;
	output wire out11_valid;
	output wire out12;
	output wire out12_valid;
	wire allDone;
	wire done12;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	wire _GEN_3 = ~emitted_4 & in0_valid;
	wire done4 = (out4_ready & _GEN_3) | emitted_4;
	reg emitted_5;
	wire _GEN_4 = ~emitted_5 & in0_valid;
	wire done5 = (out5_ready & _GEN_4) | emitted_5;
	reg emitted_6;
	wire _GEN_5 = ~emitted_6 & in0_valid;
	wire done6 = (out6_ready & _GEN_5) | emitted_6;
	reg emitted_7;
	wire _GEN_6 = ~emitted_7 & in0_valid;
	wire done7 = (out7_ready & _GEN_6) | emitted_7;
	reg emitted_8;
	wire _GEN_7 = ~emitted_8 & in0_valid;
	wire done8 = (out8_ready & _GEN_7) | emitted_8;
	reg emitted_9;
	wire _GEN_8 = ~emitted_9 & in0_valid;
	wire done9 = (out9_ready & _GEN_8) | emitted_9;
	reg emitted_10;
	wire _GEN_9 = ~emitted_10 & in0_valid;
	wire done10 = (out10_ready & _GEN_9) | emitted_10;
	reg emitted_11;
	wire _GEN_10 = ~emitted_11 & in0_valid;
	wire done11 = (out11_ready & _GEN_10) | emitted_11;
	reg emitted_12;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
			emitted_5 <= 1'h0;
			emitted_6 <= 1'h0;
			emitted_7 <= 1'h0;
			emitted_8 <= 1'h0;
			emitted_9 <= 1'h0;
			emitted_10 <= 1'h0;
			emitted_11 <= 1'h0;
			emitted_12 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
			emitted_5 <= done5 & ~allDone;
			emitted_6 <= done6 & ~allDone;
			emitted_7 <= done7 & ~allDone;
			emitted_8 <= done8 & ~allDone;
			emitted_9 <= done9 & ~allDone;
			emitted_10 <= done10 & ~allDone;
			emitted_11 <= done11 & ~allDone;
			emitted_12 <= done12 & ~allDone;
		end
	wire _GEN_11 = ~emitted_12 & in0_valid;
	assign done12 = (out12_ready & _GEN_11) | emitted_12;
	assign allDone = (((((((((((done0 & done1) & done2) & done3) & done4) & done5) & done6) & done7) & done8) & done9) & done10) & done11) & done12;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
	assign out3 = in0;
	assign out3_valid = _GEN_2;
	assign out4 = in0;
	assign out4_valid = _GEN_3;
	assign out5 = in0;
	assign out5_valid = _GEN_4;
	assign out6 = in0;
	assign out6_valid = _GEN_5;
	assign out7 = in0;
	assign out7_valid = _GEN_6;
	assign out8 = in0;
	assign out8_valid = _GEN_7;
	assign out9 = in0;
	assign out9_valid = _GEN_8;
	assign out10 = in0;
	assign out10_valid = _GEN_9;
	assign out11 = in0;
	assign out11_valid = _GEN_10;
	assign out12 = in0;
	assign out12_valid = _GEN_11;
endmodule
module handshake_fork_in_ui64_out_ui64_ui64_ui64 (
	in0,
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	in0_ready,
	out0,
	out0_valid,
	out1,
	out1_valid,
	out2,
	out2_valid
);
	input [63:0] in0;
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	output wire in0_ready;
	output wire [63:0] out0;
	output wire out0_valid;
	output wire [63:0] out1;
	output wire out1_valid;
	output wire [63:0] out2;
	output wire out2_valid;
	wire allDone;
	wire done2;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
		end
	wire _GEN_1 = ~emitted_2 & in0_valid;
	assign done2 = (out2_ready & _GEN_1) | emitted_2;
	assign allDone = (done0 & done1) & done2;
	assign in0_ready = allDone;
	assign out0 = in0;
	assign out0_valid = _GEN;
	assign out1 = in0;
	assign out1_valid = _GEN_0;
	assign out2 = in0;
	assign out2_valid = _GEN_1;
endmodule
module handshake_fork_1ins_3outs_ctrl (
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	in0_ready,
	out0_valid,
	out1_valid,
	out2_valid
);
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	output wire in0_ready;
	output wire out0_valid;
	output wire out1_valid;
	output wire out2_valid;
	wire allDone;
	wire done2;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
		end
	wire _GEN_1 = ~emitted_2 & in0_valid;
	assign done2 = (out2_ready & _GEN_1) | emitted_2;
	assign allDone = (done0 & done1) & done2;
	assign in0_ready = allDone;
	assign out0_valid = _GEN;
	assign out1_valid = _GEN_0;
	assign out2_valid = _GEN_1;
endmodule
module handshake_fork_1ins_5outs_ctrl (
	in0_valid,
	clock,
	reset,
	out0_ready,
	out1_ready,
	out2_ready,
	out3_ready,
	out4_ready,
	in0_ready,
	out0_valid,
	out1_valid,
	out2_valid,
	out3_valid,
	out4_valid
);
	input in0_valid;
	input clock;
	input reset;
	input out0_ready;
	input out1_ready;
	input out2_ready;
	input out3_ready;
	input out4_ready;
	output wire in0_ready;
	output wire out0_valid;
	output wire out1_valid;
	output wire out2_valid;
	output wire out3_valid;
	output wire out4_valid;
	wire allDone;
	wire done4;
	reg emitted_0;
	wire _GEN = ~emitted_0 & in0_valid;
	wire done0 = (out0_ready & _GEN) | emitted_0;
	reg emitted_1;
	wire _GEN_0 = ~emitted_1 & in0_valid;
	wire done1 = (out1_ready & _GEN_0) | emitted_1;
	reg emitted_2;
	wire _GEN_1 = ~emitted_2 & in0_valid;
	wire done2 = (out2_ready & _GEN_1) | emitted_2;
	reg emitted_3;
	wire _GEN_2 = ~emitted_3 & in0_valid;
	wire done3 = (out3_ready & _GEN_2) | emitted_3;
	reg emitted_4;
	always @(posedge clock)
		if (reset) begin
			emitted_0 <= 1'h0;
			emitted_1 <= 1'h0;
			emitted_2 <= 1'h0;
			emitted_3 <= 1'h0;
			emitted_4 <= 1'h0;
		end
		else begin
			emitted_0 <= done0 & ~allDone;
			emitted_1 <= done1 & ~allDone;
			emitted_2 <= done2 & ~allDone;
			emitted_3 <= done3 & ~allDone;
			emitted_4 <= done4 & ~allDone;
		end
	wire _GEN_3 = ~emitted_4 & in0_valid;
	assign done4 = (out4_ready & _GEN_3) | emitted_4;
	assign allDone = (((done0 & done1) & done2) & done3) & done4;
	assign in0_ready = allDone;
	assign out0_valid = _GEN;
	assign out1_valid = _GEN_0;
	assign out2_valid = _GEN_1;
	assign out3_valid = _GEN_2;
	assign out4_valid = _GEN_3;
endmodule
module handshake_join_3ins_1outs_ctrl (
	in0_valid,
	in1_valid,
	in2_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	in2_ready,
	out0_valid
);
	input in0_valid;
	input in1_valid;
	input in2_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire in2_ready;
	output wire out0_valid;
	wire _GEN = (in0_valid & in1_valid) & in2_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign in2_ready = _GEN_0;
	assign out0_valid = _GEN;
endmodule
module arith_addi_in_ui32_ui32_out_ui32 (
	in0,
	in0_valid,
	in1,
	in1_valid,
	out0_ready,
	in0_ready,
	in1_ready,
	out0,
	out0_valid
);
	input [31:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input out0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire [31:0] out0;
	output wire out0_valid;
	wire _GEN = in0_valid & in1_valid;
	wire _GEN_0 = out0_ready & _GEN;
	assign in0_ready = _GEN_0;
	assign in1_ready = _GEN_0;
	assign out0 = in0 + in1;
	assign out0_valid = _GEN;
endmodule
module handshake_store_in_ui64_ui32_out_ui32_ui64 (
	addrIn0,
	addrIn0_valid,
	dataIn,
	dataIn_valid,
	ctrl_valid,
	dataToMem_ready,
	addrOut0_ready,
	addrIn0_ready,
	dataIn_ready,
	ctrl_ready,
	dataToMem,
	dataToMem_valid,
	addrOut0,
	addrOut0_valid
);
	input [63:0] addrIn0;
	input addrIn0_valid;
	input [31:0] dataIn;
	input dataIn_valid;
	input ctrl_valid;
	input dataToMem_ready;
	input addrOut0_ready;
	output wire addrIn0_ready;
	output wire dataIn_ready;
	output wire ctrl_ready;
	output wire [31:0] dataToMem;
	output wire dataToMem_valid;
	output wire [63:0] addrOut0;
	output wire addrOut0_valid;
	wire _GEN = (dataIn_valid & addrIn0_valid) & ctrl_valid;
	wire _GEN_0 = (dataToMem_ready & addrOut0_ready) & _GEN;
	assign addrIn0_ready = _GEN_0;
	assign dataIn_ready = _GEN_0;
	assign ctrl_ready = _GEN_0;
	assign dataToMem = dataIn;
	assign dataToMem_valid = _GEN;
	assign addrOut0 = addrIn0;
	assign addrOut0_valid = _GEN;
endmodule
module gemm (
	in0,
	in0_valid,
	in1,
	in1_valid,
	in2_ld0_data,
	in2_ld0_data_valid,
	in3_ld0_data,
	in3_ld0_data_valid,
	in4_ld0_data,
	in4_ld0_data_valid,
	in4_st0_done_valid,
	in5_valid,
	clock,
	reset,
	out0_ready,
	in2_ld0_addr_ready,
	in3_ld0_addr_ready,
	in4_ld0_addr_ready,
	in4_st0_ready,
	in0_ready,
	in1_ready,
	in2_ld0_data_ready,
	in3_ld0_data_ready,
	in4_ld0_data_ready,
	in4_st0_done_ready,
	in5_ready,
	out0_valid,
	in2_ld0_addr,
	in2_ld0_addr_valid,
	in3_ld0_addr,
	in3_ld0_addr_valid,
	in4_ld0_addr,
	in4_ld0_addr_valid,
	in4_st0,
	in4_st0_valid
);
	input [31:0] in0;
	input in0_valid;
	input [31:0] in1;
	input in1_valid;
	input [31:0] in2_ld0_data;
	input in2_ld0_data_valid;
	input [31:0] in3_ld0_data;
	input in3_ld0_data_valid;
	input [31:0] in4_ld0_data;
	input in4_ld0_data_valid;
	input in4_st0_done_valid;
	input in5_valid;
	input clock;
	input reset;
	input out0_ready;
	input in2_ld0_addr_ready;
	input in3_ld0_addr_ready;
	input in4_ld0_addr_ready;
	input in4_st0_ready;
	output wire in0_ready;
	output wire in1_ready;
	output wire in2_ld0_data_ready;
	output wire in3_ld0_data_ready;
	output wire in4_ld0_data_ready;
	output wire in4_st0_done_ready;
	output wire in5_ready;
	output wire out0_valid;
	output wire [9:0] in2_ld0_addr;
	output wire in2_ld0_addr_valid;
	output wire [9:0] in3_ld0_addr;
	output wire in3_ld0_addr_valid;
	output wire [9:0] in4_ld0_addr;
	output wire in4_ld0_addr_valid;
	output wire [41:0] in4_st0;
	output wire in4_st0_valid;
	wire _handshake_buffer251_in0_ready;
	wire [63:0] _handshake_buffer251_out0;
	wire _handshake_buffer251_out0_valid;
	wire _arith_addi7_in0_ready;
	wire _arith_addi7_in1_ready;
	wire [63:0] _arith_addi7_out0;
	wire _arith_addi7_out0_valid;
	wire _handshake_buffer250_in0_ready;
	wire [63:0] _handshake_buffer250_out0;
	wire _handshake_buffer250_out0_valid;
	wire _arith_addi6_in0_ready;
	wire _arith_addi6_in1_ready;
	wire [63:0] _arith_addi6_out0;
	wire _arith_addi6_out0_valid;
	wire _handshake_buffer249_in0_ready;
	wire [31:0] _handshake_buffer249_out0;
	wire _handshake_buffer249_out0_valid;
	wire _handshake_buffer248_in0_ready;
	wire [63:0] _handshake_buffer248_out0;
	wire _handshake_buffer248_out0_valid;
	wire _handshake_store0_addrIn0_ready;
	wire _handshake_store0_dataIn_ready;
	wire _handshake_store0_ctrl_ready;
	wire [31:0] _handshake_store0_dataToMem;
	wire _handshake_store0_dataToMem_valid;
	wire [63:0] _handshake_store0_addrOut0;
	wire _handshake_store0_addrOut0_valid;
	wire _handshake_buffer247_in0_ready;
	wire [63:0] _handshake_buffer247_out0;
	wire _handshake_buffer247_out0_valid;
	wire _arith_addi5_in0_ready;
	wire _arith_addi5_in1_ready;
	wire [63:0] _arith_addi5_out0;
	wire _arith_addi5_out0_valid;
	wire _handshake_buffer246_in0_ready;
	wire [63:0] _handshake_buffer246_out0;
	wire _handshake_buffer246_out0_valid;
	wire _arith_muli6_in0_ready;
	wire _arith_muli6_in1_ready;
	wire [63:0] _arith_muli6_out0;
	wire _arith_muli6_out0_valid;
	wire _handshake_buffer245_in0_ready;
	wire [63:0] _handshake_buffer245_out0;
	wire _handshake_buffer245_out0_valid;
	wire _handshake_constant12_ctrl_ready;
	wire [63:0] _handshake_constant12_out0;
	wire _handshake_constant12_out0_valid;
	wire _handshake_buffer244_in0_ready;
	wire _handshake_buffer244_out0_valid;
	wire _handshake_join5_in0_ready;
	wire _handshake_join5_in1_ready;
	wire _handshake_join5_out0_valid;
	wire _handshake_buffer243_in0_ready;
	wire [63:0] _handshake_buffer243_out0;
	wire _handshake_buffer243_out0_valid;
	wire _arith_addi4_in0_ready;
	wire _arith_addi4_in1_ready;
	wire [63:0] _arith_addi4_out0;
	wire _arith_addi4_out0_valid;
	wire _handshake_buffer242_in0_ready;
	wire [31:0] _handshake_buffer242_out0;
	wire _handshake_buffer242_out0_valid;
	wire _arith_addi3_in0_ready;
	wire _arith_addi3_in1_ready;
	wire [31:0] _arith_addi3_out0;
	wire _arith_addi3_out0_valid;
	wire _handshake_buffer241_in0_ready;
	wire [31:0] _handshake_buffer241_out0;
	wire _handshake_buffer241_out0_valid;
	wire _arith_muli5_in0_ready;
	wire _arith_muli5_in1_ready;
	wire [31:0] _arith_muli5_out0;
	wire _arith_muli5_out0_valid;
	wire _handshake_buffer240_in0_ready;
	wire [31:0] _handshake_buffer240_out0;
	wire _handshake_buffer240_out0_valid;
	wire _handshake_buffer239_in0_ready;
	wire [63:0] _handshake_buffer239_out0;
	wire _handshake_buffer239_out0_valid;
	wire _handshake_load2_addrIn0_ready;
	wire _handshake_load2_dataFromMem_ready;
	wire _handshake_load2_ctrl_ready;
	wire [31:0] _handshake_load2_dataOut;
	wire _handshake_load2_dataOut_valid;
	wire [63:0] _handshake_load2_addrOut0;
	wire _handshake_load2_addrOut0_valid;
	wire _handshake_buffer238_in0_ready;
	wire [63:0] _handshake_buffer238_out0;
	wire _handshake_buffer238_out0_valid;
	wire _arith_addi2_in0_ready;
	wire _arith_addi2_in1_ready;
	wire [63:0] _arith_addi2_out0;
	wire _arith_addi2_out0_valid;
	wire _handshake_buffer237_in0_ready;
	wire [63:0] _handshake_buffer237_out0;
	wire _handshake_buffer237_out0_valid;
	wire _arith_muli4_in0_ready;
	wire _arith_muli4_in1_ready;
	wire [63:0] _arith_muli4_out0;
	wire _arith_muli4_out0_valid;
	wire _handshake_buffer236_in0_ready;
	wire [63:0] _handshake_buffer236_out0;
	wire _handshake_buffer236_out0_valid;
	wire _handshake_constant11_ctrl_ready;
	wire [63:0] _handshake_constant11_out0;
	wire _handshake_constant11_out0_valid;
	wire _handshake_buffer235_in0_ready;
	wire [31:0] _handshake_buffer235_out0;
	wire _handshake_buffer235_out0_valid;
	wire _arith_muli3_in0_ready;
	wire _arith_muli3_in1_ready;
	wire [31:0] _arith_muli3_out0;
	wire _arith_muli3_out0_valid;
	wire _handshake_buffer234_in0_ready;
	wire [31:0] _handshake_buffer234_out0;
	wire _handshake_buffer234_out0_valid;
	wire _handshake_buffer233_in0_ready;
	wire [63:0] _handshake_buffer233_out0;
	wire _handshake_buffer233_out0_valid;
	wire _handshake_load1_addrIn0_ready;
	wire _handshake_load1_dataFromMem_ready;
	wire _handshake_load1_ctrl_ready;
	wire [31:0] _handshake_load1_dataOut;
	wire _handshake_load1_dataOut_valid;
	wire [63:0] _handshake_load1_addrOut0;
	wire _handshake_load1_addrOut0_valid;
	wire _handshake_buffer232_in0_ready;
	wire [63:0] _handshake_buffer232_out0;
	wire _handshake_buffer232_out0_valid;
	wire _arith_addi1_in0_ready;
	wire _arith_addi1_in1_ready;
	wire [63:0] _arith_addi1_out0;
	wire _arith_addi1_out0_valid;
	wire _handshake_buffer231_in0_ready;
	wire [63:0] _handshake_buffer231_out0;
	wire _handshake_buffer231_out0_valid;
	wire _arith_muli2_in0_ready;
	wire _arith_muli2_in1_ready;
	wire [63:0] _arith_muli2_out0;
	wire _arith_muli2_out0_valid;
	wire _handshake_buffer230_in0_ready;
	wire [63:0] _handshake_buffer230_out0;
	wire _handshake_buffer230_out0_valid;
	wire _handshake_constant10_ctrl_ready;
	wire [63:0] _handshake_constant10_out0;
	wire _handshake_constant10_out0_valid;
	wire _handshake_buffer229_in0_ready;
	wire _handshake_buffer229_out0_valid;
	wire _handshake_join4_in0_ready;
	wire _handshake_join4_in1_ready;
	wire _handshake_join4_in2_ready;
	wire _handshake_join4_out0_valid;
	wire _handshake_buffer228_in0_ready;
	wire _handshake_buffer228_out0_valid;
	wire _handshake_buffer227_in0_ready;
	wire _handshake_buffer227_out0_valid;
	wire _handshake_buffer226_in0_ready;
	wire _handshake_buffer226_out0_valid;
	wire _handshake_buffer225_in0_ready;
	wire _handshake_buffer225_out0_valid;
	wire _handshake_buffer224_in0_ready;
	wire _handshake_buffer224_out0_valid;
	wire _handshake_fork31_in0_ready;
	wire _handshake_fork31_out0_valid;
	wire _handshake_fork31_out1_valid;
	wire _handshake_fork31_out2_valid;
	wire _handshake_fork31_out3_valid;
	wire _handshake_fork31_out4_valid;
	wire _handshake_buffer223_in0_ready;
	wire _handshake_buffer223_out0_valid;
	wire _handshake_buffer222_in0_ready;
	wire _handshake_buffer222_out0_valid;
	wire _handshake_buffer221_in0_ready;
	wire _handshake_buffer221_out0_valid;
	wire _handshake_fork30_in0_ready;
	wire _handshake_fork30_out0_valid;
	wire _handshake_fork30_out1_valid;
	wire _handshake_fork30_out2_valid;
	wire _handshake_buffer220_in0_ready;
	wire _handshake_buffer220_out0_valid;
	wire _handshake_buffer219_in0_ready;
	wire _handshake_buffer219_out0_valid;
	wire _handshake_cond_br27_cond_ready;
	wire _handshake_cond_br27_data_ready;
	wire _handshake_cond_br27_outTrue_valid;
	wire _handshake_cond_br27_outFalse_valid;
	wire _handshake_buffer218_in0_ready;
	wire [63:0] _handshake_buffer218_out0;
	wire _handshake_buffer218_out0_valid;
	wire _handshake_buffer217_in0_ready;
	wire [63:0] _handshake_buffer217_out0;
	wire _handshake_buffer217_out0_valid;
	wire _handshake_fork29_in0_ready;
	wire [63:0] _handshake_fork29_out0;
	wire _handshake_fork29_out0_valid;
	wire [63:0] _handshake_fork29_out1;
	wire _handshake_fork29_out1_valid;
	wire _handshake_sink10_in0_ready;
	wire _handshake_buffer216_in0_ready;
	wire [63:0] _handshake_buffer216_out0;
	wire _handshake_buffer216_out0_valid;
	wire _handshake_cond_br26_cond_ready;
	wire _handshake_cond_br26_data_ready;
	wire [63:0] _handshake_cond_br26_outTrue;
	wire _handshake_cond_br26_outTrue_valid;
	wire [63:0] _handshake_cond_br26_outFalse;
	wire _handshake_cond_br26_outFalse_valid;
	wire _handshake_sink9_in0_ready;
	wire _handshake_buffer215_in0_ready;
	wire [63:0] _handshake_buffer215_out0;
	wire _handshake_buffer215_out0_valid;
	wire _handshake_cond_br25_cond_ready;
	wire _handshake_cond_br25_data_ready;
	wire [63:0] _handshake_cond_br25_outTrue;
	wire _handshake_cond_br25_outTrue_valid;
	wire [63:0] _handshake_cond_br25_outFalse;
	wire _handshake_cond_br25_outFalse_valid;
	wire _handshake_buffer214_in0_ready;
	wire [63:0] _handshake_buffer214_out0;
	wire _handshake_buffer214_out0_valid;
	wire _handshake_buffer213_in0_ready;
	wire [63:0] _handshake_buffer213_out0;
	wire _handshake_buffer213_out0_valid;
	wire _handshake_fork28_in0_ready;
	wire [63:0] _handshake_fork28_out0;
	wire _handshake_fork28_out0_valid;
	wire [63:0] _handshake_fork28_out1;
	wire _handshake_fork28_out1_valid;
	wire _handshake_buffer212_in0_ready;
	wire [63:0] _handshake_buffer212_out0;
	wire _handshake_buffer212_out0_valid;
	wire _handshake_buffer211_in0_ready;
	wire [63:0] _handshake_buffer211_out0;
	wire _handshake_buffer211_out0_valid;
	wire _handshake_fork27_in0_ready;
	wire [63:0] _handshake_fork27_out0;
	wire _handshake_fork27_out0_valid;
	wire [63:0] _handshake_fork27_out1;
	wire _handshake_fork27_out1_valid;
	wire _handshake_buffer210_in0_ready;
	wire [63:0] _handshake_buffer210_out0;
	wire _handshake_buffer210_out0_valid;
	wire _handshake_buffer209_in0_ready;
	wire [63:0] _handshake_buffer209_out0;
	wire _handshake_buffer209_out0_valid;
	wire _handshake_cond_br24_cond_ready;
	wire _handshake_cond_br24_data_ready;
	wire [63:0] _handshake_cond_br24_outTrue;
	wire _handshake_cond_br24_outTrue_valid;
	wire [63:0] _handshake_cond_br24_outFalse;
	wire _handshake_cond_br24_outFalse_valid;
	wire _handshake_buffer208_in0_ready;
	wire [63:0] _handshake_buffer208_out0;
	wire _handshake_buffer208_out0_valid;
	wire _handshake_buffer207_in0_ready;
	wire [63:0] _handshake_buffer207_out0;
	wire _handshake_buffer207_out0_valid;
	wire _handshake_fork26_in0_ready;
	wire [63:0] _handshake_fork26_out0;
	wire _handshake_fork26_out0_valid;
	wire [63:0] _handshake_fork26_out1;
	wire _handshake_fork26_out1_valid;
	wire _handshake_buffer206_in0_ready;
	wire [63:0] _handshake_buffer206_out0;
	wire _handshake_buffer206_out0_valid;
	wire _handshake_buffer205_in0_ready;
	wire [63:0] _handshake_buffer205_out0;
	wire _handshake_buffer205_out0_valid;
	wire _handshake_cond_br23_cond_ready;
	wire _handshake_cond_br23_data_ready;
	wire [63:0] _handshake_cond_br23_outTrue;
	wire _handshake_cond_br23_outTrue_valid;
	wire [63:0] _handshake_cond_br23_outFalse;
	wire _handshake_cond_br23_outFalse_valid;
	wire _handshake_buffer204_in0_ready;
	wire [63:0] _handshake_buffer204_out0;
	wire _handshake_buffer204_out0_valid;
	wire _handshake_buffer203_in0_ready;
	wire [63:0] _handshake_buffer203_out0;
	wire _handshake_buffer203_out0_valid;
	wire _handshake_cond_br22_cond_ready;
	wire _handshake_cond_br22_data_ready;
	wire [63:0] _handshake_cond_br22_outTrue;
	wire _handshake_cond_br22_outTrue_valid;
	wire [63:0] _handshake_cond_br22_outFalse;
	wire _handshake_cond_br22_outFalse_valid;
	wire _handshake_buffer202_in0_ready;
	wire [63:0] _handshake_buffer202_out0;
	wire _handshake_buffer202_out0_valid;
	wire _handshake_buffer201_in0_ready;
	wire [63:0] _handshake_buffer201_out0;
	wire _handshake_buffer201_out0_valid;
	wire _handshake_fork25_in0_ready;
	wire [63:0] _handshake_fork25_out0;
	wire _handshake_fork25_out0_valid;
	wire [63:0] _handshake_fork25_out1;
	wire _handshake_fork25_out1_valid;
	wire _handshake_buffer200_in0_ready;
	wire [63:0] _handshake_buffer200_out0;
	wire _handshake_buffer200_out0_valid;
	wire _handshake_buffer199_in0_ready;
	wire [63:0] _handshake_buffer199_out0;
	wire _handshake_buffer199_out0_valid;
	wire _handshake_fork24_in0_ready;
	wire [63:0] _handshake_fork24_out0;
	wire _handshake_fork24_out0_valid;
	wire [63:0] _handshake_fork24_out1;
	wire _handshake_fork24_out1_valid;
	wire _handshake_buffer198_in0_ready;
	wire [63:0] _handshake_buffer198_out0;
	wire _handshake_buffer198_out0_valid;
	wire _handshake_buffer197_in0_ready;
	wire [63:0] _handshake_buffer197_out0;
	wire _handshake_buffer197_out0_valid;
	wire _handshake_cond_br21_cond_ready;
	wire _handshake_cond_br21_data_ready;
	wire [63:0] _handshake_cond_br21_outTrue;
	wire _handshake_cond_br21_outTrue_valid;
	wire [63:0] _handshake_cond_br21_outFalse;
	wire _handshake_cond_br21_outFalse_valid;
	wire _handshake_buffer196_in0_ready;
	wire [63:0] _handshake_buffer196_out0;
	wire _handshake_buffer196_out0_valid;
	wire _handshake_buffer195_in0_ready;
	wire [63:0] _handshake_buffer195_out0;
	wire _handshake_buffer195_out0_valid;
	wire _handshake_cond_br20_cond_ready;
	wire _handshake_cond_br20_data_ready;
	wire [63:0] _handshake_cond_br20_outTrue;
	wire _handshake_cond_br20_outTrue_valid;
	wire [63:0] _handshake_cond_br20_outFalse;
	wire _handshake_cond_br20_outFalse_valid;
	wire _handshake_buffer194_in0_ready;
	wire [63:0] _handshake_buffer194_out0;
	wire _handshake_buffer194_out0_valid;
	wire _handshake_buffer193_in0_ready;
	wire [63:0] _handshake_buffer193_out0;
	wire _handshake_buffer193_out0_valid;
	wire _handshake_cond_br19_cond_ready;
	wire _handshake_cond_br19_data_ready;
	wire [63:0] _handshake_cond_br19_outTrue;
	wire _handshake_cond_br19_outTrue_valid;
	wire [63:0] _handshake_cond_br19_outFalse;
	wire _handshake_cond_br19_outFalse_valid;
	wire _handshake_buffer192_in0_ready;
	wire [31:0] _handshake_buffer192_out0;
	wire _handshake_buffer192_out0_valid;
	wire _handshake_buffer191_in0_ready;
	wire [31:0] _handshake_buffer191_out0;
	wire _handshake_buffer191_out0_valid;
	wire _handshake_cond_br18_cond_ready;
	wire _handshake_cond_br18_data_ready;
	wire [31:0] _handshake_cond_br18_outTrue;
	wire _handshake_cond_br18_outTrue_valid;
	wire [31:0] _handshake_cond_br18_outFalse;
	wire _handshake_cond_br18_outFalse_valid;
	wire _handshake_buffer190_in0_ready;
	wire [31:0] _handshake_buffer190_out0;
	wire _handshake_buffer190_out0_valid;
	wire _handshake_buffer189_in0_ready;
	wire [31:0] _handshake_buffer189_out0;
	wire _handshake_buffer189_out0_valid;
	wire _handshake_fork23_in0_ready;
	wire [31:0] _handshake_fork23_out0;
	wire _handshake_fork23_out0_valid;
	wire [31:0] _handshake_fork23_out1;
	wire _handshake_fork23_out1_valid;
	wire _handshake_buffer188_in0_ready;
	wire [31:0] _handshake_buffer188_out0;
	wire _handshake_buffer188_out0_valid;
	wire _handshake_buffer187_in0_ready;
	wire [31:0] _handshake_buffer187_out0;
	wire _handshake_buffer187_out0_valid;
	wire _handshake_cond_br17_cond_ready;
	wire _handshake_cond_br17_data_ready;
	wire [31:0] _handshake_cond_br17_outTrue;
	wire _handshake_cond_br17_outTrue_valid;
	wire [31:0] _handshake_cond_br17_outFalse;
	wire _handshake_cond_br17_outFalse_valid;
	wire _handshake_buffer186_in0_ready;
	wire [31:0] _handshake_buffer186_out0;
	wire _handshake_buffer186_out0_valid;
	wire _handshake_buffer185_in0_ready;
	wire [31:0] _handshake_buffer185_out0;
	wire _handshake_buffer185_out0_valid;
	wire _handshake_cond_br16_cond_ready;
	wire _handshake_cond_br16_data_ready;
	wire [31:0] _handshake_cond_br16_outTrue;
	wire _handshake_cond_br16_outTrue_valid;
	wire [31:0] _handshake_cond_br16_outFalse;
	wire _handshake_cond_br16_outFalse_valid;
	wire _handshake_buffer184_in0_ready;
	wire [63:0] _handshake_buffer184_out0;
	wire _handshake_buffer184_out0_valid;
	wire _handshake_buffer183_in0_ready;
	wire [63:0] _handshake_buffer183_out0;
	wire _handshake_buffer183_out0_valid;
	wire _handshake_buffer182_in0_ready;
	wire [63:0] _handshake_buffer182_out0;
	wire _handshake_buffer182_out0_valid;
	wire _handshake_fork22_in0_ready;
	wire [63:0] _handshake_fork22_out0;
	wire _handshake_fork22_out0_valid;
	wire [63:0] _handshake_fork22_out1;
	wire _handshake_fork22_out1_valid;
	wire [63:0] _handshake_fork22_out2;
	wire _handshake_fork22_out2_valid;
	wire _handshake_sink8_in0_ready;
	wire _handshake_buffer181_in0_ready;
	wire [63:0] _handshake_buffer181_out0;
	wire _handshake_buffer181_out0_valid;
	wire _handshake_cond_br15_cond_ready;
	wire _handshake_cond_br15_data_ready;
	wire [63:0] _handshake_cond_br15_outTrue;
	wire _handshake_cond_br15_outTrue_valid;
	wire [63:0] _handshake_cond_br15_outFalse;
	wire _handshake_cond_br15_outFalse_valid;
	wire _handshake_buffer180_in0_ready;
	wire _handshake_buffer180_out0;
	wire _handshake_buffer180_out0_valid;
	wire _handshake_buffer179_in0_ready;
	wire _handshake_buffer179_out0;
	wire _handshake_buffer179_out0_valid;
	wire _handshake_buffer178_in0_ready;
	wire _handshake_buffer178_out0;
	wire _handshake_buffer178_out0_valid;
	wire _handshake_buffer177_in0_ready;
	wire _handshake_buffer177_out0;
	wire _handshake_buffer177_out0_valid;
	wire _handshake_buffer176_in0_ready;
	wire _handshake_buffer176_out0;
	wire _handshake_buffer176_out0_valid;
	wire _handshake_buffer175_in0_ready;
	wire _handshake_buffer175_out0;
	wire _handshake_buffer175_out0_valid;
	wire _handshake_buffer174_in0_ready;
	wire _handshake_buffer174_out0;
	wire _handshake_buffer174_out0_valid;
	wire _handshake_buffer173_in0_ready;
	wire _handshake_buffer173_out0;
	wire _handshake_buffer173_out0_valid;
	wire _handshake_buffer172_in0_ready;
	wire _handshake_buffer172_out0;
	wire _handshake_buffer172_out0_valid;
	wire _handshake_buffer171_in0_ready;
	wire _handshake_buffer171_out0;
	wire _handshake_buffer171_out0_valid;
	wire _handshake_buffer170_in0_ready;
	wire _handshake_buffer170_out0;
	wire _handshake_buffer170_out0_valid;
	wire _handshake_buffer169_in0_ready;
	wire _handshake_buffer169_out0;
	wire _handshake_buffer169_out0_valid;
	wire _handshake_buffer168_in0_ready;
	wire _handshake_buffer168_out0;
	wire _handshake_buffer168_out0_valid;
	wire _handshake_fork21_in0_ready;
	wire _handshake_fork21_out0;
	wire _handshake_fork21_out0_valid;
	wire _handshake_fork21_out1;
	wire _handshake_fork21_out1_valid;
	wire _handshake_fork21_out2;
	wire _handshake_fork21_out2_valid;
	wire _handshake_fork21_out3;
	wire _handshake_fork21_out3_valid;
	wire _handshake_fork21_out4;
	wire _handshake_fork21_out4_valid;
	wire _handshake_fork21_out5;
	wire _handshake_fork21_out5_valid;
	wire _handshake_fork21_out6;
	wire _handshake_fork21_out6_valid;
	wire _handshake_fork21_out7;
	wire _handshake_fork21_out7_valid;
	wire _handshake_fork21_out8;
	wire _handshake_fork21_out8_valid;
	wire _handshake_fork21_out9;
	wire _handshake_fork21_out9_valid;
	wire _handshake_fork21_out10;
	wire _handshake_fork21_out10_valid;
	wire _handshake_fork21_out11;
	wire _handshake_fork21_out11_valid;
	wire _handshake_fork21_out12;
	wire _handshake_fork21_out12_valid;
	wire _handshake_buffer167_in0_ready;
	wire _handshake_buffer167_out0;
	wire _handshake_buffer167_out0_valid;
	wire _arith_cmpi2_in0_ready;
	wire _arith_cmpi2_in1_ready;
	wire _arith_cmpi2_out0;
	wire _arith_cmpi2_out0_valid;
	wire _handshake_buffer166_in0_ready;
	wire [63:0] _handshake_buffer166_out0;
	wire _handshake_buffer166_out0_valid;
	wire _handshake_buffer165_in0_ready;
	wire [63:0] _handshake_buffer165_out0;
	wire _handshake_buffer165_out0_valid;
	wire _handshake_buffer164_in0_ready;
	wire [63:0] _handshake_buffer164_out0;
	wire _handshake_buffer164_out0_valid;
	wire _handshake_buffer163_in0_ready;
	wire [63:0] _handshake_buffer163_out0;
	wire _handshake_buffer163_out0_valid;
	wire _handshake_buffer162_in0_ready;
	wire [63:0] _handshake_buffer162_out0;
	wire _handshake_buffer162_out0_valid;
	wire _handshake_buffer161_in0_ready;
	wire [63:0] _handshake_buffer161_out0;
	wire _handshake_buffer161_out0_valid;
	wire _handshake_buffer160_in0_ready;
	wire [63:0] _handshake_buffer160_out0;
	wire _handshake_buffer160_out0_valid;
	wire _handshake_buffer159_in0_ready;
	wire [63:0] _handshake_buffer159_out0;
	wire _handshake_buffer159_out0_valid;
	wire _handshake_buffer158_in0_ready;
	wire [63:0] _handshake_buffer158_out0;
	wire _handshake_buffer158_out0_valid;
	wire _handshake_buffer157_in0_ready;
	wire [63:0] _handshake_buffer157_out0;
	wire _handshake_buffer157_out0_valid;
	wire _handshake_buffer156_in0_ready;
	wire [63:0] _handshake_buffer156_out0;
	wire _handshake_buffer156_out0_valid;
	wire _handshake_buffer155_in0_ready;
	wire [63:0] _handshake_buffer155_out0;
	wire _handshake_buffer155_out0_valid;
	wire _handshake_fork20_in0_ready;
	wire [63:0] _handshake_fork20_out0;
	wire _handshake_fork20_out0_valid;
	wire [63:0] _handshake_fork20_out1;
	wire _handshake_fork20_out1_valid;
	wire [63:0] _handshake_fork20_out2;
	wire _handshake_fork20_out2_valid;
	wire [63:0] _handshake_fork20_out3;
	wire _handshake_fork20_out3_valid;
	wire [63:0] _handshake_fork20_out4;
	wire _handshake_fork20_out4_valid;
	wire [63:0] _handshake_fork20_out5;
	wire _handshake_fork20_out5_valid;
	wire [63:0] _handshake_fork20_out6;
	wire _handshake_fork20_out6_valid;
	wire [63:0] _handshake_fork20_out7;
	wire _handshake_fork20_out7_valid;
	wire [63:0] _handshake_fork20_out8;
	wire _handshake_fork20_out8_valid;
	wire [63:0] _handshake_fork20_out9;
	wire _handshake_fork20_out9_valid;
	wire [63:0] _handshake_fork20_out10;
	wire _handshake_fork20_out10_valid;
	wire [63:0] _handshake_fork20_out11;
	wire _handshake_fork20_out11_valid;
	wire _handshake_buffer154_in0_ready;
	wire _handshake_buffer154_out0_valid;
	wire _handshake_buffer153_in0_ready;
	wire [63:0] _handshake_buffer153_out0;
	wire _handshake_buffer153_out0_valid;
	wire _handshake_control_merge1_in0_ready;
	wire _handshake_control_merge1_in1_ready;
	wire _handshake_control_merge1_dataOut_valid;
	wire [63:0] _handshake_control_merge1_index;
	wire _handshake_control_merge1_index_valid;
	wire _handshake_buffer152_in0_ready;
	wire [63:0] _handshake_buffer152_out0;
	wire _handshake_buffer152_out0_valid;
	wire _handshake_mux25_select_ready;
	wire _handshake_mux25_in0_ready;
	wire _handshake_mux25_in1_ready;
	wire [63:0] _handshake_mux25_out0;
	wire _handshake_mux25_out0_valid;
	wire _handshake_buffer151_in0_ready;
	wire [63:0] _handshake_buffer151_out0;
	wire _handshake_buffer151_out0_valid;
	wire _handshake_buffer150_in0_ready;
	wire [63:0] _handshake_buffer150_out0;
	wire _handshake_buffer150_out0_valid;
	wire _handshake_fork19_in0_ready;
	wire [63:0] _handshake_fork19_out0;
	wire _handshake_fork19_out0_valid;
	wire [63:0] _handshake_fork19_out1;
	wire _handshake_fork19_out1_valid;
	wire _handshake_buffer149_in0_ready;
	wire [63:0] _handshake_buffer149_out0;
	wire _handshake_buffer149_out0_valid;
	wire _handshake_mux24_select_ready;
	wire _handshake_mux24_in0_ready;
	wire _handshake_mux24_in1_ready;
	wire [63:0] _handshake_mux24_out0;
	wire _handshake_mux24_out0_valid;
	wire _handshake_buffer148_in0_ready;
	wire [63:0] _handshake_buffer148_out0;
	wire _handshake_buffer148_out0_valid;
	wire _handshake_mux23_select_ready;
	wire _handshake_mux23_in0_ready;
	wire _handshake_mux23_in1_ready;
	wire [63:0] _handshake_mux23_out0;
	wire _handshake_mux23_out0_valid;
	wire _handshake_buffer147_in0_ready;
	wire [63:0] _handshake_buffer147_out0;
	wire _handshake_buffer147_out0_valid;
	wire _handshake_mux22_select_ready;
	wire _handshake_mux22_in0_ready;
	wire _handshake_mux22_in1_ready;
	wire [63:0] _handshake_mux22_out0;
	wire _handshake_mux22_out0_valid;
	wire _handshake_buffer146_in0_ready;
	wire [63:0] _handshake_buffer146_out0;
	wire _handshake_buffer146_out0_valid;
	wire _handshake_mux21_select_ready;
	wire _handshake_mux21_in0_ready;
	wire _handshake_mux21_in1_ready;
	wire [63:0] _handshake_mux21_out0;
	wire _handshake_mux21_out0_valid;
	wire _handshake_buffer145_in0_ready;
	wire [63:0] _handshake_buffer145_out0;
	wire _handshake_buffer145_out0_valid;
	wire _handshake_mux20_select_ready;
	wire _handshake_mux20_in0_ready;
	wire _handshake_mux20_in1_ready;
	wire [63:0] _handshake_mux20_out0;
	wire _handshake_mux20_out0_valid;
	wire _handshake_buffer144_in0_ready;
	wire [63:0] _handshake_buffer144_out0;
	wire _handshake_buffer144_out0_valid;
	wire _handshake_mux19_select_ready;
	wire _handshake_mux19_in0_ready;
	wire _handshake_mux19_in1_ready;
	wire [63:0] _handshake_mux19_out0;
	wire _handshake_mux19_out0_valid;
	wire _handshake_buffer143_in0_ready;
	wire [63:0] _handshake_buffer143_out0;
	wire _handshake_buffer143_out0_valid;
	wire _handshake_mux18_select_ready;
	wire _handshake_mux18_in0_ready;
	wire _handshake_mux18_in1_ready;
	wire [63:0] _handshake_mux18_out0;
	wire _handshake_mux18_out0_valid;
	wire _handshake_buffer142_in0_ready;
	wire [31:0] _handshake_buffer142_out0;
	wire _handshake_buffer142_out0_valid;
	wire _handshake_mux17_select_ready;
	wire _handshake_mux17_in0_ready;
	wire _handshake_mux17_in1_ready;
	wire [31:0] _handshake_mux17_out0;
	wire _handshake_mux17_out0_valid;
	wire _handshake_buffer141_in0_ready;
	wire [31:0] _handshake_buffer141_out0;
	wire _handshake_buffer141_out0_valid;
	wire _handshake_mux16_select_ready;
	wire _handshake_mux16_in0_ready;
	wire _handshake_mux16_in1_ready;
	wire [31:0] _handshake_mux16_out0;
	wire _handshake_mux16_out0_valid;
	wire _handshake_buffer140_in0_ready;
	wire [31:0] _handshake_buffer140_out0;
	wire _handshake_buffer140_out0_valid;
	wire _handshake_mux15_select_ready;
	wire _handshake_mux15_in0_ready;
	wire _handshake_mux15_in1_ready;
	wire [31:0] _handshake_mux15_out0;
	wire _handshake_mux15_out0_valid;
	wire _handshake_buffer139_in0_ready;
	wire [63:0] _handshake_buffer139_out0;
	wire _handshake_buffer139_out0_valid;
	wire _handshake_buffer138_in0_ready;
	wire [63:0] _handshake_buffer138_out0;
	wire _handshake_buffer138_out0_valid;
	wire _handshake_fork18_in0_ready;
	wire [63:0] _handshake_fork18_out0;
	wire _handshake_fork18_out0_valid;
	wire [63:0] _handshake_fork18_out1;
	wire _handshake_fork18_out1_valid;
	wire _handshake_buffer137_in0_ready;
	wire [63:0] _handshake_buffer137_out0;
	wire _handshake_buffer137_out0_valid;
	wire _handshake_mux14_select_ready;
	wire _handshake_mux14_in0_ready;
	wire _handshake_mux14_in1_ready;
	wire [63:0] _handshake_mux14_out0;
	wire _handshake_mux14_out0_valid;
	wire _handshake_buffer136_in0_ready;
	wire [63:0] _handshake_buffer136_out0;
	wire _handshake_buffer136_out0_valid;
	wire _handshake_constant9_ctrl_ready;
	wire [63:0] _handshake_constant9_out0;
	wire _handshake_constant9_out0_valid;
	wire _handshake_buffer135_in0_ready;
	wire [63:0] _handshake_buffer135_out0;
	wire _handshake_buffer135_out0_valid;
	wire _handshake_constant8_ctrl_ready;
	wire [63:0] _handshake_constant8_out0;
	wire _handshake_constant8_out0_valid;
	wire _handshake_buffer134_in0_ready;
	wire [63:0] _handshake_buffer134_out0;
	wire _handshake_buffer134_out0_valid;
	wire _handshake_constant7_ctrl_ready;
	wire [63:0] _handshake_constant7_out0;
	wire _handshake_constant7_out0_valid;
	wire _handshake_buffer133_in0_ready;
	wire [31:0] _handshake_buffer133_out0;
	wire _handshake_buffer133_out0_valid;
	wire _arith_muli1_in0_ready;
	wire _arith_muli1_in1_ready;
	wire [31:0] _arith_muli1_out0;
	wire _arith_muli1_out0_valid;
	wire _handshake_buffer132_in0_ready;
	wire [31:0] _handshake_buffer132_out0;
	wire _handshake_buffer132_out0_valid;
	wire _handshake_buffer131_in0_ready;
	wire [63:0] _handshake_buffer131_out0;
	wire _handshake_buffer131_out0_valid;
	wire _handshake_load0_addrIn0_ready;
	wire _handshake_load0_dataFromMem_ready;
	wire _handshake_load0_ctrl_ready;
	wire [31:0] _handshake_load0_dataOut;
	wire _handshake_load0_dataOut_valid;
	wire [63:0] _handshake_load0_addrOut0;
	wire _handshake_load0_addrOut0_valid;
	wire _handshake_buffer130_in0_ready;
	wire [63:0] _handshake_buffer130_out0;
	wire _handshake_buffer130_out0_valid;
	wire _arith_addi0_in0_ready;
	wire _arith_addi0_in1_ready;
	wire [63:0] _arith_addi0_out0;
	wire _arith_addi0_out0_valid;
	wire _handshake_buffer129_in0_ready;
	wire [63:0] _handshake_buffer129_out0;
	wire _handshake_buffer129_out0_valid;
	wire _arith_muli0_in0_ready;
	wire _arith_muli0_in1_ready;
	wire [63:0] _arith_muli0_out0;
	wire _arith_muli0_out0_valid;
	wire _handshake_buffer128_in0_ready;
	wire [63:0] _handshake_buffer128_out0;
	wire _handshake_buffer128_out0_valid;
	wire _handshake_constant6_ctrl_ready;
	wire [63:0] _handshake_constant6_out0;
	wire _handshake_constant6_out0_valid;
	wire _handshake_buffer127_in0_ready;
	wire _handshake_buffer127_out0_valid;
	wire _handshake_join3_in0_ready;
	wire _handshake_join3_in1_ready;
	wire _handshake_join3_out0_valid;
	wire _handshake_buffer126_in0_ready;
	wire _handshake_buffer126_out0_valid;
	wire _handshake_buffer125_in0_ready;
	wire _handshake_buffer125_out0_valid;
	wire _handshake_buffer124_in0_ready;
	wire _handshake_buffer124_out0_valid;
	wire _handshake_buffer123_in0_ready;
	wire _handshake_buffer123_out0_valid;
	wire _handshake_buffer122_in0_ready;
	wire _handshake_buffer122_out0_valid;
	wire _handshake_buffer121_in0_ready;
	wire _handshake_buffer121_out0_valid;
	wire _handshake_fork17_in0_ready;
	wire _handshake_fork17_out0_valid;
	wire _handshake_fork17_out1_valid;
	wire _handshake_fork17_out2_valid;
	wire _handshake_fork17_out3_valid;
	wire _handshake_fork17_out4_valid;
	wire _handshake_fork17_out5_valid;
	wire _handshake_buffer120_in0_ready;
	wire _handshake_buffer120_out0_valid;
	wire _handshake_buffer119_in0_ready;
	wire _handshake_buffer119_out0_valid;
	wire _handshake_cond_br14_cond_ready;
	wire _handshake_cond_br14_data_ready;
	wire _handshake_cond_br14_outTrue_valid;
	wire _handshake_cond_br14_outFalse_valid;
	wire _handshake_sink7_in0_ready;
	wire _handshake_buffer118_in0_ready;
	wire [63:0] _handshake_buffer118_out0;
	wire _handshake_buffer118_out0_valid;
	wire _handshake_cond_br13_cond_ready;
	wire _handshake_cond_br13_data_ready;
	wire [63:0] _handshake_cond_br13_outTrue;
	wire _handshake_cond_br13_outTrue_valid;
	wire [63:0] _handshake_cond_br13_outFalse;
	wire _handshake_cond_br13_outFalse_valid;
	wire _handshake_sink6_in0_ready;
	wire _handshake_buffer117_in0_ready;
	wire [63:0] _handshake_buffer117_out0;
	wire _handshake_buffer117_out0_valid;
	wire _handshake_cond_br12_cond_ready;
	wire _handshake_cond_br12_data_ready;
	wire [63:0] _handshake_cond_br12_outTrue;
	wire _handshake_cond_br12_outTrue_valid;
	wire [63:0] _handshake_cond_br12_outFalse;
	wire _handshake_cond_br12_outFalse_valid;
	wire _handshake_buffer116_in0_ready;
	wire [63:0] _handshake_buffer116_out0;
	wire _handshake_buffer116_out0_valid;
	wire _handshake_buffer115_in0_ready;
	wire [63:0] _handshake_buffer115_out0;
	wire _handshake_buffer115_out0_valid;
	wire _handshake_fork16_in0_ready;
	wire [63:0] _handshake_fork16_out0;
	wire _handshake_fork16_out0_valid;
	wire [63:0] _handshake_fork16_out1;
	wire _handshake_fork16_out1_valid;
	wire _handshake_buffer114_in0_ready;
	wire [63:0] _handshake_buffer114_out0;
	wire _handshake_buffer114_out0_valid;
	wire _handshake_buffer113_in0_ready;
	wire [63:0] _handshake_buffer113_out0;
	wire _handshake_buffer113_out0_valid;
	wire _handshake_cond_br11_cond_ready;
	wire _handshake_cond_br11_data_ready;
	wire [63:0] _handshake_cond_br11_outTrue;
	wire _handshake_cond_br11_outTrue_valid;
	wire [63:0] _handshake_cond_br11_outFalse;
	wire _handshake_cond_br11_outFalse_valid;
	wire _handshake_buffer112_in0_ready;
	wire [63:0] _handshake_buffer112_out0;
	wire _handshake_buffer112_out0_valid;
	wire _handshake_buffer111_in0_ready;
	wire [63:0] _handshake_buffer111_out0;
	wire _handshake_buffer111_out0_valid;
	wire _handshake_fork15_in0_ready;
	wire [63:0] _handshake_fork15_out0;
	wire _handshake_fork15_out0_valid;
	wire [63:0] _handshake_fork15_out1;
	wire _handshake_fork15_out1_valid;
	wire _handshake_buffer110_in0_ready;
	wire [63:0] _handshake_buffer110_out0;
	wire _handshake_buffer110_out0_valid;
	wire _handshake_buffer109_in0_ready;
	wire [63:0] _handshake_buffer109_out0;
	wire _handshake_buffer109_out0_valid;
	wire _handshake_cond_br10_cond_ready;
	wire _handshake_cond_br10_data_ready;
	wire [63:0] _handshake_cond_br10_outTrue;
	wire _handshake_cond_br10_outTrue_valid;
	wire [63:0] _handshake_cond_br10_outFalse;
	wire _handshake_cond_br10_outFalse_valid;
	wire _handshake_buffer108_in0_ready;
	wire [63:0] _handshake_buffer108_out0;
	wire _handshake_buffer108_out0_valid;
	wire _handshake_buffer107_in0_ready;
	wire [63:0] _handshake_buffer107_out0;
	wire _handshake_buffer107_out0_valid;
	wire _handshake_cond_br9_cond_ready;
	wire _handshake_cond_br9_data_ready;
	wire [63:0] _handshake_cond_br9_outTrue;
	wire _handshake_cond_br9_outTrue_valid;
	wire [63:0] _handshake_cond_br9_outFalse;
	wire _handshake_cond_br9_outFalse_valid;
	wire _handshake_buffer106_in0_ready;
	wire [31:0] _handshake_buffer106_out0;
	wire _handshake_buffer106_out0_valid;
	wire _handshake_buffer105_in0_ready;
	wire [31:0] _handshake_buffer105_out0;
	wire _handshake_buffer105_out0_valid;
	wire _handshake_fork14_in0_ready;
	wire [31:0] _handshake_fork14_out0;
	wire _handshake_fork14_out0_valid;
	wire [31:0] _handshake_fork14_out1;
	wire _handshake_fork14_out1_valid;
	wire _handshake_buffer104_in0_ready;
	wire [31:0] _handshake_buffer104_out0;
	wire _handshake_buffer104_out0_valid;
	wire _handshake_buffer103_in0_ready;
	wire [31:0] _handshake_buffer103_out0;
	wire _handshake_buffer103_out0_valid;
	wire _handshake_cond_br8_cond_ready;
	wire _handshake_cond_br8_data_ready;
	wire [31:0] _handshake_cond_br8_outTrue;
	wire _handshake_cond_br8_outTrue_valid;
	wire [31:0] _handshake_cond_br8_outFalse;
	wire _handshake_cond_br8_outFalse_valid;
	wire _handshake_buffer102_in0_ready;
	wire [31:0] _handshake_buffer102_out0;
	wire _handshake_buffer102_out0_valid;
	wire _handshake_buffer101_in0_ready;
	wire [31:0] _handshake_buffer101_out0;
	wire _handshake_buffer101_out0_valid;
	wire _handshake_cond_br7_cond_ready;
	wire _handshake_cond_br7_data_ready;
	wire [31:0] _handshake_cond_br7_outTrue;
	wire _handshake_cond_br7_outTrue_valid;
	wire [31:0] _handshake_cond_br7_outFalse;
	wire _handshake_cond_br7_outFalse_valid;
	wire _handshake_buffer100_in0_ready;
	wire [63:0] _handshake_buffer100_out0;
	wire _handshake_buffer100_out0_valid;
	wire _handshake_buffer99_in0_ready;
	wire [63:0] _handshake_buffer99_out0;
	wire _handshake_buffer99_out0_valid;
	wire _handshake_fork13_in0_ready;
	wire [63:0] _handshake_fork13_out0;
	wire _handshake_fork13_out0_valid;
	wire [63:0] _handshake_fork13_out1;
	wire _handshake_fork13_out1_valid;
	wire _handshake_sink5_in0_ready;
	wire _handshake_buffer98_in0_ready;
	wire [63:0] _handshake_buffer98_out0;
	wire _handshake_buffer98_out0_valid;
	wire _handshake_cond_br6_cond_ready;
	wire _handshake_cond_br6_data_ready;
	wire [63:0] _handshake_cond_br6_outTrue;
	wire _handshake_cond_br6_outTrue_valid;
	wire [63:0] _handshake_cond_br6_outFalse;
	wire _handshake_cond_br6_outFalse_valid;
	wire _handshake_buffer97_in0_ready;
	wire _handshake_buffer97_out0;
	wire _handshake_buffer97_out0_valid;
	wire _handshake_buffer96_in0_ready;
	wire _handshake_buffer96_out0;
	wire _handshake_buffer96_out0_valid;
	wire _handshake_buffer95_in0_ready;
	wire _handshake_buffer95_out0;
	wire _handshake_buffer95_out0_valid;
	wire _handshake_buffer94_in0_ready;
	wire _handshake_buffer94_out0;
	wire _handshake_buffer94_out0_valid;
	wire _handshake_buffer93_in0_ready;
	wire _handshake_buffer93_out0;
	wire _handshake_buffer93_out0_valid;
	wire _handshake_buffer92_in0_ready;
	wire _handshake_buffer92_out0;
	wire _handshake_buffer92_out0_valid;
	wire _handshake_buffer91_in0_ready;
	wire _handshake_buffer91_out0;
	wire _handshake_buffer91_out0_valid;
	wire _handshake_buffer90_in0_ready;
	wire _handshake_buffer90_out0;
	wire _handshake_buffer90_out0_valid;
	wire _handshake_buffer89_in0_ready;
	wire _handshake_buffer89_out0;
	wire _handshake_buffer89_out0_valid;
	wire _handshake_fork12_in0_ready;
	wire _handshake_fork12_out0;
	wire _handshake_fork12_out0_valid;
	wire _handshake_fork12_out1;
	wire _handshake_fork12_out1_valid;
	wire _handshake_fork12_out2;
	wire _handshake_fork12_out2_valid;
	wire _handshake_fork12_out3;
	wire _handshake_fork12_out3_valid;
	wire _handshake_fork12_out4;
	wire _handshake_fork12_out4_valid;
	wire _handshake_fork12_out5;
	wire _handshake_fork12_out5_valid;
	wire _handshake_fork12_out6;
	wire _handshake_fork12_out6_valid;
	wire _handshake_fork12_out7;
	wire _handshake_fork12_out7_valid;
	wire _handshake_fork12_out8;
	wire _handshake_fork12_out8_valid;
	wire _handshake_buffer88_in0_ready;
	wire _handshake_buffer88_out0;
	wire _handshake_buffer88_out0_valid;
	wire _arith_cmpi1_in0_ready;
	wire _arith_cmpi1_in1_ready;
	wire _arith_cmpi1_out0;
	wire _arith_cmpi1_out0_valid;
	wire _handshake_buffer87_in0_ready;
	wire [63:0] _handshake_buffer87_out0;
	wire _handshake_buffer87_out0_valid;
	wire _handshake_buffer86_in0_ready;
	wire [63:0] _handshake_buffer86_out0;
	wire _handshake_buffer86_out0_valid;
	wire _handshake_buffer85_in0_ready;
	wire [63:0] _handshake_buffer85_out0;
	wire _handshake_buffer85_out0_valid;
	wire _handshake_buffer84_in0_ready;
	wire [63:0] _handshake_buffer84_out0;
	wire _handshake_buffer84_out0_valid;
	wire _handshake_buffer83_in0_ready;
	wire [63:0] _handshake_buffer83_out0;
	wire _handshake_buffer83_out0_valid;
	wire _handshake_buffer82_in0_ready;
	wire [63:0] _handshake_buffer82_out0;
	wire _handshake_buffer82_out0_valid;
	wire _handshake_buffer81_in0_ready;
	wire [63:0] _handshake_buffer81_out0;
	wire _handshake_buffer81_out0_valid;
	wire _handshake_buffer80_in0_ready;
	wire [63:0] _handshake_buffer80_out0;
	wire _handshake_buffer80_out0_valid;
	wire _handshake_fork11_in0_ready;
	wire [63:0] _handshake_fork11_out0;
	wire _handshake_fork11_out0_valid;
	wire [63:0] _handshake_fork11_out1;
	wire _handshake_fork11_out1_valid;
	wire [63:0] _handshake_fork11_out2;
	wire _handshake_fork11_out2_valid;
	wire [63:0] _handshake_fork11_out3;
	wire _handshake_fork11_out3_valid;
	wire [63:0] _handshake_fork11_out4;
	wire _handshake_fork11_out4_valid;
	wire [63:0] _handshake_fork11_out5;
	wire _handshake_fork11_out5_valid;
	wire [63:0] _handshake_fork11_out6;
	wire _handshake_fork11_out6_valid;
	wire [63:0] _handshake_fork11_out7;
	wire _handshake_fork11_out7_valid;
	wire _handshake_buffer79_in0_ready;
	wire _handshake_buffer79_out0_valid;
	wire _handshake_buffer78_in0_ready;
	wire [63:0] _handshake_buffer78_out0;
	wire _handshake_buffer78_out0_valid;
	wire _handshake_control_merge0_in0_ready;
	wire _handshake_control_merge0_in1_ready;
	wire _handshake_control_merge0_dataOut_valid;
	wire [63:0] _handshake_control_merge0_index;
	wire _handshake_control_merge0_index_valid;
	wire _handshake_buffer77_in0_ready;
	wire [63:0] _handshake_buffer77_out0;
	wire _handshake_buffer77_out0_valid;
	wire _handshake_mux13_select_ready;
	wire _handshake_mux13_in0_ready;
	wire _handshake_mux13_in1_ready;
	wire [63:0] _handshake_mux13_out0;
	wire _handshake_mux13_out0_valid;
	wire _handshake_buffer76_in0_ready;
	wire [63:0] _handshake_buffer76_out0;
	wire _handshake_buffer76_out0_valid;
	wire _handshake_buffer75_in0_ready;
	wire [63:0] _handshake_buffer75_out0;
	wire _handshake_buffer75_out0_valid;
	wire _handshake_fork10_in0_ready;
	wire [63:0] _handshake_fork10_out0;
	wire _handshake_fork10_out0_valid;
	wire [63:0] _handshake_fork10_out1;
	wire _handshake_fork10_out1_valid;
	wire _handshake_buffer74_in0_ready;
	wire [63:0] _handshake_buffer74_out0;
	wire _handshake_buffer74_out0_valid;
	wire _handshake_mux12_select_ready;
	wire _handshake_mux12_in0_ready;
	wire _handshake_mux12_in1_ready;
	wire [63:0] _handshake_mux12_out0;
	wire _handshake_mux12_out0_valid;
	wire _handshake_buffer73_in0_ready;
	wire [63:0] _handshake_buffer73_out0;
	wire _handshake_buffer73_out0_valid;
	wire _handshake_mux11_select_ready;
	wire _handshake_mux11_in0_ready;
	wire _handshake_mux11_in1_ready;
	wire [63:0] _handshake_mux11_out0;
	wire _handshake_mux11_out0_valid;
	wire _handshake_buffer72_in0_ready;
	wire [63:0] _handshake_buffer72_out0;
	wire _handshake_buffer72_out0_valid;
	wire _handshake_mux10_select_ready;
	wire _handshake_mux10_in0_ready;
	wire _handshake_mux10_in1_ready;
	wire [63:0] _handshake_mux10_out0;
	wire _handshake_mux10_out0_valid;
	wire _handshake_buffer71_in0_ready;
	wire [63:0] _handshake_buffer71_out0;
	wire _handshake_buffer71_out0_valid;
	wire _handshake_mux9_select_ready;
	wire _handshake_mux9_in0_ready;
	wire _handshake_mux9_in1_ready;
	wire [63:0] _handshake_mux9_out0;
	wire _handshake_mux9_out0_valid;
	wire _handshake_buffer70_in0_ready;
	wire [31:0] _handshake_buffer70_out0;
	wire _handshake_buffer70_out0_valid;
	wire _handshake_mux8_select_ready;
	wire _handshake_mux8_in0_ready;
	wire _handshake_mux8_in1_ready;
	wire [31:0] _handshake_mux8_out0;
	wire _handshake_mux8_out0_valid;
	wire _handshake_buffer69_in0_ready;
	wire [31:0] _handshake_buffer69_out0;
	wire _handshake_buffer69_out0_valid;
	wire _handshake_mux7_select_ready;
	wire _handshake_mux7_in0_ready;
	wire _handshake_mux7_in1_ready;
	wire [31:0] _handshake_mux7_out0;
	wire _handshake_mux7_out0_valid;
	wire _handshake_buffer68_in0_ready;
	wire [63:0] _handshake_buffer68_out0;
	wire _handshake_buffer68_out0_valid;
	wire _handshake_buffer67_in0_ready;
	wire [63:0] _handshake_buffer67_out0;
	wire _handshake_buffer67_out0_valid;
	wire _handshake_fork9_in0_ready;
	wire [63:0] _handshake_fork9_out0;
	wire _handshake_fork9_out0_valid;
	wire [63:0] _handshake_fork9_out1;
	wire _handshake_fork9_out1_valid;
	wire _handshake_buffer66_in0_ready;
	wire [63:0] _handshake_buffer66_out0;
	wire _handshake_buffer66_out0_valid;
	wire _handshake_mux6_select_ready;
	wire _handshake_mux6_in0_ready;
	wire _handshake_mux6_in1_ready;
	wire [63:0] _handshake_mux6_out0;
	wire _handshake_mux6_out0_valid;
	wire _handshake_buffer65_in0_ready;
	wire [63:0] _handshake_buffer65_out0;
	wire _handshake_buffer65_out0_valid;
	wire _handshake_constant5_ctrl_ready;
	wire [63:0] _handshake_constant5_out0;
	wire _handshake_constant5_out0_valid;
	wire _handshake_buffer64_in0_ready;
	wire [63:0] _handshake_buffer64_out0;
	wire _handshake_buffer64_out0_valid;
	wire _handshake_constant4_ctrl_ready;
	wire [63:0] _handshake_constant4_out0;
	wire _handshake_constant4_out0_valid;
	wire _handshake_buffer63_in0_ready;
	wire [63:0] _handshake_buffer63_out0;
	wire _handshake_buffer63_out0_valid;
	wire _handshake_constant3_ctrl_ready;
	wire [63:0] _handshake_constant3_out0;
	wire _handshake_constant3_out0_valid;
	wire _handshake_buffer62_in0_ready;
	wire _handshake_buffer62_out0_valid;
	wire _handshake_buffer61_in0_ready;
	wire _handshake_buffer61_out0_valid;
	wire _handshake_buffer60_in0_ready;
	wire _handshake_buffer60_out0_valid;
	wire _handshake_buffer59_in0_ready;
	wire _handshake_buffer59_out0_valid;
	wire _handshake_fork8_in0_ready;
	wire _handshake_fork8_out0_valid;
	wire _handshake_fork8_out1_valid;
	wire _handshake_fork8_out2_valid;
	wire _handshake_fork8_out3_valid;
	wire _handshake_buffer58_in0_ready;
	wire _handshake_buffer58_out0_valid;
	wire _handshake_buffer57_in0_ready;
	wire _handshake_cond_br5_cond_ready;
	wire _handshake_cond_br5_data_ready;
	wire _handshake_cond_br5_outTrue_valid;
	wire _handshake_cond_br5_outFalse_valid;
	wire _handshake_sink4_in0_ready;
	wire _handshake_buffer56_in0_ready;
	wire [63:0] _handshake_buffer56_out0;
	wire _handshake_buffer56_out0_valid;
	wire _handshake_cond_br4_cond_ready;
	wire _handshake_cond_br4_data_ready;
	wire [63:0] _handshake_cond_br4_outTrue;
	wire _handshake_cond_br4_outTrue_valid;
	wire [63:0] _handshake_cond_br4_outFalse;
	wire _handshake_cond_br4_outFalse_valid;
	wire _handshake_sink3_in0_ready;
	wire _handshake_buffer55_in0_ready;
	wire [63:0] _handshake_buffer55_out0;
	wire _handshake_buffer55_out0_valid;
	wire _handshake_cond_br3_cond_ready;
	wire _handshake_cond_br3_data_ready;
	wire [63:0] _handshake_cond_br3_outTrue;
	wire _handshake_cond_br3_outTrue_valid;
	wire [63:0] _handshake_cond_br3_outFalse;
	wire _handshake_cond_br3_outFalse_valid;
	wire _handshake_sink2_in0_ready;
	wire _handshake_buffer54_in0_ready;
	wire [31:0] _handshake_buffer54_out0;
	wire _handshake_buffer54_out0_valid;
	wire _handshake_cond_br2_cond_ready;
	wire _handshake_cond_br2_data_ready;
	wire [31:0] _handshake_cond_br2_outTrue;
	wire _handshake_cond_br2_outTrue_valid;
	wire [31:0] _handshake_cond_br2_outFalse;
	wire _handshake_cond_br2_outFalse_valid;
	wire _handshake_sink1_in0_ready;
	wire _handshake_buffer53_in0_ready;
	wire [31:0] _handshake_buffer53_out0;
	wire _handshake_buffer53_out0_valid;
	wire _handshake_cond_br1_cond_ready;
	wire _handshake_cond_br1_data_ready;
	wire [31:0] _handshake_cond_br1_outTrue;
	wire _handshake_cond_br1_outTrue_valid;
	wire [31:0] _handshake_cond_br1_outFalse;
	wire _handshake_cond_br1_outFalse_valid;
	wire _handshake_sink0_in0_ready;
	wire _handshake_buffer52_in0_ready;
	wire [63:0] _handshake_buffer52_out0;
	wire _handshake_buffer52_out0_valid;
	wire _handshake_cond_br0_cond_ready;
	wire _handshake_cond_br0_data_ready;
	wire [63:0] _handshake_cond_br0_outTrue;
	wire _handshake_cond_br0_outTrue_valid;
	wire [63:0] _handshake_cond_br0_outFalse;
	wire _handshake_cond_br0_outFalse_valid;
	wire _handshake_buffer51_in0_ready;
	wire _handshake_buffer51_out0;
	wire _handshake_buffer51_out0_valid;
	wire _handshake_buffer50_in0_ready;
	wire _handshake_buffer50_out0;
	wire _handshake_buffer50_out0_valid;
	wire _handshake_buffer49_in0_ready;
	wire _handshake_buffer49_out0;
	wire _handshake_buffer49_out0_valid;
	wire _handshake_buffer48_in0_ready;
	wire _handshake_buffer48_out0;
	wire _handshake_buffer48_out0_valid;
	wire _handshake_buffer47_in0_ready;
	wire _handshake_buffer47_out0;
	wire _handshake_buffer47_out0_valid;
	wire _handshake_buffer46_in0_ready;
	wire _handshake_buffer46_out0;
	wire _handshake_buffer46_out0_valid;
	wire _handshake_fork7_in0_ready;
	wire _handshake_fork7_out0;
	wire _handshake_fork7_out0_valid;
	wire _handshake_fork7_out1;
	wire _handshake_fork7_out1_valid;
	wire _handshake_fork7_out2;
	wire _handshake_fork7_out2_valid;
	wire _handshake_fork7_out3;
	wire _handshake_fork7_out3_valid;
	wire _handshake_fork7_out4;
	wire _handshake_fork7_out4_valid;
	wire _handshake_fork7_out5;
	wire _handshake_fork7_out5_valid;
	wire _handshake_fork7_out6;
	wire _handshake_fork7_out6_valid;
	wire _handshake_buffer45_in0_ready;
	wire _handshake_buffer45_out0;
	wire _handshake_buffer45_out0_valid;
	wire _arith_cmpi0_in0_ready;
	wire _arith_cmpi0_in1_ready;
	wire _arith_cmpi0_out0;
	wire _arith_cmpi0_out0_valid;
	wire _handshake_buffer44_in0_ready;
	wire [63:0] _handshake_buffer44_out0;
	wire _handshake_buffer44_out0_valid;
	wire _handshake_mux5_select_ready;
	wire _handshake_mux5_in0_ready;
	wire _handshake_mux5_in1_ready;
	wire [63:0] _handshake_mux5_out0;
	wire _handshake_mux5_out0_valid;
	wire _handshake_buffer43_in0_ready;
	wire [63:0] _handshake_buffer43_out0;
	wire _handshake_buffer43_out0_valid;
	wire _handshake_buffer42_in0_ready;
	wire [63:0] _handshake_buffer42_out0;
	wire _handshake_buffer42_out0_valid;
	wire _handshake_fork6_in0_ready;
	wire [63:0] _handshake_fork6_out0;
	wire _handshake_fork6_out0_valid;
	wire [63:0] _handshake_fork6_out1;
	wire _handshake_fork6_out1_valid;
	wire _handshake_buffer41_in0_ready;
	wire [63:0] _handshake_buffer41_out0;
	wire _handshake_buffer41_out0_valid;
	wire _handshake_mux4_select_ready;
	wire _handshake_mux4_in0_ready;
	wire _handshake_mux4_in1_ready;
	wire [63:0] _handshake_mux4_out0;
	wire _handshake_mux4_out0_valid;
	wire _handshake_buffer40_in0_ready;
	wire [31:0] _handshake_buffer40_out0;
	wire _handshake_buffer40_out0_valid;
	wire _handshake_mux3_select_ready;
	wire _handshake_mux3_in0_ready;
	wire _handshake_mux3_in1_ready;
	wire [31:0] _handshake_mux3_out0;
	wire _handshake_mux3_out0_valid;
	wire _handshake_buffer39_in0_ready;
	wire [31:0] _handshake_buffer39_out0;
	wire _handshake_buffer39_out0_valid;
	wire _handshake_mux2_select_ready;
	wire _handshake_mux2_in0_ready;
	wire _handshake_mux2_in1_ready;
	wire [31:0] _handshake_mux2_out0;
	wire _handshake_mux2_out0_valid;
	wire _handshake_buffer38_in0_ready;
	wire [63:0] _handshake_buffer38_out0;
	wire _handshake_buffer38_out0_valid;
	wire _handshake_buffer37_in0_ready;
	wire [63:0] _handshake_buffer37_out0;
	wire _handshake_buffer37_out0_valid;
	wire _handshake_fork5_in0_ready;
	wire [63:0] _handshake_fork5_out0;
	wire _handshake_fork5_out0_valid;
	wire [63:0] _handshake_fork5_out1;
	wire _handshake_fork5_out1_valid;
	wire _handshake_buffer36_in0_ready;
	wire [63:0] _handshake_buffer36_out0;
	wire _handshake_buffer36_out0_valid;
	wire _handshake_mux1_select_ready;
	wire _handshake_mux1_in0_ready;
	wire _handshake_mux1_in1_ready;
	wire [63:0] _handshake_mux1_out0;
	wire _handshake_mux1_out0_valid;
	wire _handshake_buffer35_in0_ready;
	wire _handshake_buffer35_out0_valid;
	wire _handshake_mux0_select_ready;
	wire _handshake_mux0_in0_ready;
	wire _handshake_mux0_in1_ready;
	wire _handshake_mux0_out0_valid;
	wire _handshake_buffer34_in0_ready;
	wire _handshake_buffer34_out0;
	wire _handshake_buffer34_out0_valid;
	wire _handshake_buffer33_in0_ready;
	wire _handshake_buffer33_out0;
	wire _handshake_buffer33_out0_valid;
	wire _handshake_buffer32_in0_ready;
	wire _handshake_buffer32_out0;
	wire _handshake_buffer32_out0_valid;
	wire _handshake_buffer31_in0_ready;
	wire _handshake_buffer31_out0;
	wire _handshake_buffer31_out0_valid;
	wire _handshake_buffer30_in0_ready;
	wire _handshake_buffer30_out0;
	wire _handshake_buffer30_out0_valid;
	wire _handshake_buffer29_in0_ready;
	wire _handshake_buffer29_out0;
	wire _handshake_buffer29_out0_valid;
	wire _handshake_fork4_in0_ready;
	wire _handshake_fork4_out0;
	wire _handshake_fork4_out0_valid;
	wire _handshake_fork4_out1;
	wire _handshake_fork4_out1_valid;
	wire _handshake_fork4_out2;
	wire _handshake_fork4_out2_valid;
	wire _handshake_fork4_out3;
	wire _handshake_fork4_out3_valid;
	wire _handshake_fork4_out4;
	wire _handshake_fork4_out4_valid;
	wire _handshake_fork4_out5;
	wire _handshake_fork4_out5_valid;
	wire _handshake_buffer28_in0_ready;
	wire _handshake_buffer28_out0;
	wire _handshake_buffer28_out0_valid;
	wire _handshake_buffer27_in0_ready;
	wire [63:0] _handshake_buffer27_out0;
	wire _handshake_buffer27_out0_valid;
	wire _handshake_constant2_ctrl_ready;
	wire [63:0] _handshake_constant2_out0;
	wire _handshake_constant2_out0_valid;
	wire _handshake_buffer26_in0_ready;
	wire [63:0] _handshake_buffer26_out0;
	wire _handshake_buffer26_out0_valid;
	wire _handshake_constant1_ctrl_ready;
	wire [63:0] _handshake_constant1_out0;
	wire _handshake_constant1_out0_valid;
	wire _handshake_buffer25_in0_ready;
	wire [63:0] _handshake_buffer25_out0;
	wire _handshake_buffer25_out0_valid;
	wire _handshake_constant0_ctrl_ready;
	wire [63:0] _handshake_constant0_out0;
	wire _handshake_constant0_out0_valid;
	wire _handshake_buffer24_in0_ready;
	wire _arith_index_cast3_in0_ready;
	wire [9:0] _arith_index_cast3_out0;
	wire _arith_index_cast3_out0_valid;
	wire _handshake_buffer23_in0_ready;
	wire _handshake_buffer23_out0_valid;
	wire _handshake_join2_in0_ready;
	wire _handshake_join2_out0_valid;
	wire _handshake_buffer22_in0_ready;
	wire [31:0] _handshake_buffer22_out0;
	wire _handshake_buffer22_out0_valid;
	wire _handshake_buffer21_in0_ready;
	wire [31:0] _handshake_buffer21_out0;
	wire _handshake_buffer21_out0_valid;
	wire _handshake_fork3_in0_ready;
	wire [31:0] _handshake_fork3_out0;
	wire _handshake_fork3_out0_valid;
	wire [31:0] _handshake_fork3_out1;
	wire _handshake_fork3_out1_valid;
	wire _handshake_buffer20_in0_ready;
	wire _arith_index_cast2_in0_ready;
	wire [9:0] _arith_index_cast2_out0;
	wire _arith_index_cast2_out0_valid;
	wire _handshake_buffer19_in0_ready;
	wire _handshake_buffer19_out0_valid;
	wire _handshake_join1_in0_ready;
	wire _handshake_join1_out0_valid;
	wire _handshake_buffer18_in0_ready;
	wire [31:0] _handshake_buffer18_out0;
	wire _handshake_buffer18_out0_valid;
	wire _handshake_buffer17_in0_ready;
	wire [31:0] _handshake_buffer17_out0;
	wire _handshake_buffer17_out0_valid;
	wire _handshake_fork2_in0_ready;
	wire [31:0] _handshake_fork2_out0;
	wire _handshake_fork2_out0_valid;
	wire [31:0] _handshake_fork2_out1;
	wire _handshake_fork2_out1_valid;
	wire _handshake_buffer16_in0_ready;
	wire _hw_struct_create0_in0_ready;
	wire _hw_struct_create0_in1_ready;
	wire [41:0] _hw_struct_create0_out0;
	wire _hw_struct_create0_out0_valid;
	wire _handshake_buffer15_in0_ready;
	wire [9:0] _handshake_buffer15_out0;
	wire _handshake_buffer15_out0_valid;
	wire _arith_index_cast1_in0_ready;
	wire [9:0] _arith_index_cast1_out0;
	wire _arith_index_cast1_out0_valid;
	wire _handshake_buffer14_in0_ready;
	wire _arith_index_cast0_in0_ready;
	wire [9:0] _arith_index_cast0_out0;
	wire _arith_index_cast0_out0_valid;
	wire _handshake_buffer13_in0_ready;
	wire _handshake_buffer13_out0_valid;
	wire _handshake_join0_in0_ready;
	wire _handshake_join0_out0_valid;
	wire _handshake_buffer12_in0_ready;
	wire [31:0] _handshake_buffer12_out0;
	wire _handshake_buffer12_out0_valid;
	wire _handshake_buffer11_in0_ready;
	wire [31:0] _handshake_buffer11_out0;
	wire _handshake_buffer11_out0_valid;
	wire _handshake_fork1_in0_ready;
	wire [31:0] _handshake_fork1_out0;
	wire _handshake_fork1_out0_valid;
	wire [31:0] _handshake_fork1_out1;
	wire _handshake_fork1_out1_valid;
	wire _handshake_buffer10_in0_ready;
	wire _handshake_buffer10_out0_valid;
	wire _handshake_buffer9_in0_ready;
	wire _handshake_buffer9_out0_valid;
	wire _handshake_buffer8_in0_ready;
	wire _handshake_buffer8_out0_valid;
	wire _handshake_buffer7_in0_ready;
	wire _handshake_buffer7_out0_valid;
	wire _handshake_fork0_in0_ready;
	wire _handshake_fork0_out0_valid;
	wire _handshake_fork0_out1_valid;
	wire _handshake_fork0_out2_valid;
	wire _handshake_fork0_out3_valid;
	wire [31:0] _handshake_buffer6_out0;
	wire _handshake_buffer6_out0_valid;
	wire [31:0] _handshake_buffer5_out0;
	wire _handshake_buffer5_out0_valid;
	wire [31:0] _handshake_buffer4_out0;
	wire _handshake_buffer4_out0_valid;
	wire [31:0] _handshake_buffer3_out0;
	wire _handshake_buffer3_out0_valid;
	wire [31:0] _handshake_buffer2_out0;
	wire _handshake_buffer2_out0_valid;
	wire _handshake_buffer1_out0_valid;
	wire _handshake_buffer0_out0_valid;
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer0(
		.in0_valid(in5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork0_in0_ready),
		.in0_ready(in5_ready),
		.out0_valid(_handshake_buffer0_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer1(
		.in0_valid(in4_st0_done_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join5_in1_ready),
		.in0_ready(in4_st0_done_ready),
		.out0_valid(_handshake_buffer1_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer2(
		.in0(in4_ld0_data),
		.in0_valid(in4_ld0_data_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork1_in0_ready),
		.in0_ready(in4_ld0_data_ready),
		.out0(_handshake_buffer2_out0),
		.out0_valid(_handshake_buffer2_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer3(
		.in0(in3_ld0_data),
		.in0_valid(in3_ld0_data_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork2_in0_ready),
		.in0_ready(in3_ld0_data_ready),
		.out0(_handshake_buffer3_out0),
		.out0_valid(_handshake_buffer3_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer4(
		.in0(in2_ld0_data),
		.in0_valid(in2_ld0_data_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork3_in0_ready),
		.in0_ready(in2_ld0_data_ready),
		.out0(_handshake_buffer4_out0),
		.out0_valid(_handshake_buffer4_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer5(
		.in0(in1),
		.in0_valid(in1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux3_in0_ready),
		.in0_ready(in1_ready),
		.out0(_handshake_buffer5_out0),
		.out0_valid(_handshake_buffer5_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer6(
		.in0(in0),
		.in0_valid(in0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux2_in0_ready),
		.in0_ready(in0_ready),
		.out0(_handshake_buffer6_out0),
		.out0_valid(_handshake_buffer6_out0_valid)
	);
	handshake_fork_1ins_4outs_ctrl handshake_fork0(
		.in0_valid(_handshake_buffer0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer10_in0_ready),
		.out1_ready(_handshake_buffer9_in0_ready),
		.out2_ready(_handshake_buffer8_in0_ready),
		.out3_ready(_handshake_buffer7_in0_ready),
		.in0_ready(_handshake_fork0_in0_ready),
		.out0_valid(_handshake_fork0_out0_valid),
		.out1_valid(_handshake_fork0_out1_valid),
		.out2_valid(_handshake_fork0_out2_valid),
		.out3_valid(_handshake_fork0_out3_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer7(
		.in0_valid(_handshake_fork0_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant2_ctrl_ready),
		.in0_ready(_handshake_buffer7_in0_ready),
		.out0_valid(_handshake_buffer7_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer8(
		.in0_valid(_handshake_fork0_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant1_ctrl_ready),
		.in0_ready(_handshake_buffer8_in0_ready),
		.out0_valid(_handshake_buffer8_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer9(
		.in0_valid(_handshake_fork0_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant0_ctrl_ready),
		.in0_ready(_handshake_buffer9_in0_ready),
		.out0_valid(_handshake_buffer9_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer10(
		.in0_valid(_handshake_fork0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux0_in0_ready),
		.in0_ready(_handshake_buffer10_in0_ready),
		.out0_valid(_handshake_buffer10_out0_valid)
	);
	handshake_fork_in_ui32_out_ui32_ui32 handshake_fork1(
		.in0(_handshake_buffer2_out0),
		.in0_valid(_handshake_buffer2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer12_in0_ready),
		.out1_ready(_handshake_buffer11_in0_ready),
		.in0_ready(_handshake_fork1_in0_ready),
		.out0(_handshake_fork1_out0),
		.out0_valid(_handshake_fork1_out0_valid),
		.out1(_handshake_fork1_out1),
		.out1_valid(_handshake_fork1_out1_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer11(
		.in0(_handshake_fork1_out1),
		.in0_valid(_handshake_fork1_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join0_in0_ready),
		.in0_ready(_handshake_buffer11_in0_ready),
		.out0(_handshake_buffer11_out0),
		.out0_valid(_handshake_buffer11_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer12(
		.in0(_handshake_fork1_out0),
		.in0_valid(_handshake_fork1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load0_dataFromMem_ready),
		.in0_ready(_handshake_buffer12_in0_ready),
		.out0(_handshake_buffer12_out0),
		.out0_valid(_handshake_buffer12_out0_valid)
	);
	handshake_join_in_ui32_1ins_1outs_ctrl handshake_join0(
		.in0(_handshake_buffer11_out0),
		.in0_valid(_handshake_buffer11_out0_valid),
		.out0_ready(_handshake_buffer13_in0_ready),
		.in0_ready(_handshake_join0_in0_ready),
		.out0_valid(_handshake_join0_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer13(
		.in0_valid(_handshake_join0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join3_in1_ready),
		.in0_ready(_handshake_buffer13_in0_ready),
		.out0_valid(_handshake_buffer13_out0_valid)
	);
	arith_index_cast_in_ui64_out_ui10 arith_index_cast0(
		.in0(_handshake_buffer131_out0),
		.in0_valid(_handshake_buffer131_out0_valid),
		.out0_ready(_handshake_buffer14_in0_ready),
		.in0_ready(_arith_index_cast0_in0_ready),
		.out0(_arith_index_cast0_out0),
		.out0_valid(_arith_index_cast0_out0_valid)
	);
	handshake_buffer_in_ui10_out_ui10_2slots_seq handshake_buffer14(
		.in0(_arith_index_cast0_out0),
		.in0_valid(_arith_index_cast0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(in4_ld0_addr_ready),
		.in0_ready(_handshake_buffer14_in0_ready),
		.out0(in4_ld0_addr),
		.out0_valid(in4_ld0_addr_valid)
	);
	arith_index_cast_in_ui64_out_ui10 arith_index_cast1(
		.in0(_handshake_buffer248_out0),
		.in0_valid(_handshake_buffer248_out0_valid),
		.out0_ready(_handshake_buffer15_in0_ready),
		.in0_ready(_arith_index_cast1_in0_ready),
		.out0(_arith_index_cast1_out0),
		.out0_valid(_arith_index_cast1_out0_valid)
	);
	handshake_buffer_in_ui10_out_ui10_2slots_seq handshake_buffer15(
		.in0(_arith_index_cast1_out0),
		.in0_valid(_arith_index_cast1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_hw_struct_create0_in0_ready),
		.in0_ready(_handshake_buffer15_in0_ready),
		.out0(_handshake_buffer15_out0),
		.out0_valid(_handshake_buffer15_out0_valid)
	);
	hw_struct_create_in_ui10_ui32_out_struct_address_ui10_data_ui32 hw_struct_create0(
		.in0(_handshake_buffer15_out0),
		.in0_valid(_handshake_buffer15_out0_valid),
		.in1(_handshake_buffer249_out0),
		.in1_valid(_handshake_buffer249_out0_valid),
		.out0_ready(_handshake_buffer16_in0_ready),
		.in0_ready(_hw_struct_create0_in0_ready),
		.in1_ready(_hw_struct_create0_in1_ready),
		.out0(_hw_struct_create0_out0),
		.out0_valid(_hw_struct_create0_out0_valid)
	);
	handshake_buffer_in_struct_address_ui10_data_ui32_out_struct_address_ui10_data_ui32_2slots_seq handshake_buffer16(
		.in0(_hw_struct_create0_out0),
		.in0_valid(_hw_struct_create0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(in4_st0_ready),
		.in0_ready(_handshake_buffer16_in0_ready),
		.out0(in4_st0),
		.out0_valid(in4_st0_valid)
	);
	handshake_fork_in_ui32_out_ui32_ui32 handshake_fork2(
		.in0(_handshake_buffer3_out0),
		.in0_valid(_handshake_buffer3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer18_in0_ready),
		.out1_ready(_handshake_buffer17_in0_ready),
		.in0_ready(_handshake_fork2_in0_ready),
		.out0(_handshake_fork2_out0),
		.out0_valid(_handshake_fork2_out0_valid),
		.out1(_handshake_fork2_out1),
		.out1_valid(_handshake_fork2_out1_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer17(
		.in0(_handshake_fork2_out1),
		.in0_valid(_handshake_fork2_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join1_in0_ready),
		.in0_ready(_handshake_buffer17_in0_ready),
		.out0(_handshake_buffer17_out0),
		.out0_valid(_handshake_buffer17_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer18(
		.in0(_handshake_fork2_out0),
		.in0_valid(_handshake_fork2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load2_dataFromMem_ready),
		.in0_ready(_handshake_buffer18_in0_ready),
		.out0(_handshake_buffer18_out0),
		.out0_valid(_handshake_buffer18_out0_valid)
	);
	handshake_join_in_ui32_1ins_1outs_ctrl handshake_join1(
		.in0(_handshake_buffer17_out0),
		.in0_valid(_handshake_buffer17_out0_valid),
		.out0_ready(_handshake_buffer19_in0_ready),
		.in0_ready(_handshake_join1_in0_ready),
		.out0_valid(_handshake_join1_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer19(
		.in0_valid(_handshake_join1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join4_in2_ready),
		.in0_ready(_handshake_buffer19_in0_ready),
		.out0_valid(_handshake_buffer19_out0_valid)
	);
	arith_index_cast_in_ui64_out_ui10 arith_index_cast2(
		.in0(_handshake_buffer239_out0),
		.in0_valid(_handshake_buffer239_out0_valid),
		.out0_ready(_handshake_buffer20_in0_ready),
		.in0_ready(_arith_index_cast2_in0_ready),
		.out0(_arith_index_cast2_out0),
		.out0_valid(_arith_index_cast2_out0_valid)
	);
	handshake_buffer_in_ui10_out_ui10_2slots_seq handshake_buffer20(
		.in0(_arith_index_cast2_out0),
		.in0_valid(_arith_index_cast2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(in3_ld0_addr_ready),
		.in0_ready(_handshake_buffer20_in0_ready),
		.out0(in3_ld0_addr),
		.out0_valid(in3_ld0_addr_valid)
	);
	handshake_fork_in_ui32_out_ui32_ui32 handshake_fork3(
		.in0(_handshake_buffer4_out0),
		.in0_valid(_handshake_buffer4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer22_in0_ready),
		.out1_ready(_handshake_buffer21_in0_ready),
		.in0_ready(_handshake_fork3_in0_ready),
		.out0(_handshake_fork3_out0),
		.out0_valid(_handshake_fork3_out0_valid),
		.out1(_handshake_fork3_out1),
		.out1_valid(_handshake_fork3_out1_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer21(
		.in0(_handshake_fork3_out1),
		.in0_valid(_handshake_fork3_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join2_in0_ready),
		.in0_ready(_handshake_buffer21_in0_ready),
		.out0(_handshake_buffer21_out0),
		.out0_valid(_handshake_buffer21_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer22(
		.in0(_handshake_fork3_out0),
		.in0_valid(_handshake_fork3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load1_dataFromMem_ready),
		.in0_ready(_handshake_buffer22_in0_ready),
		.out0(_handshake_buffer22_out0),
		.out0_valid(_handshake_buffer22_out0_valid)
	);
	handshake_join_in_ui32_1ins_1outs_ctrl handshake_join2(
		.in0(_handshake_buffer21_out0),
		.in0_valid(_handshake_buffer21_out0_valid),
		.out0_ready(_handshake_buffer23_in0_ready),
		.in0_ready(_handshake_join2_in0_ready),
		.out0_valid(_handshake_join2_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer23(
		.in0_valid(_handshake_join2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join4_in1_ready),
		.in0_ready(_handshake_buffer23_in0_ready),
		.out0_valid(_handshake_buffer23_out0_valid)
	);
	arith_index_cast_in_ui64_out_ui10 arith_index_cast3(
		.in0(_handshake_buffer233_out0),
		.in0_valid(_handshake_buffer233_out0_valid),
		.out0_ready(_handshake_buffer24_in0_ready),
		.in0_ready(_arith_index_cast3_in0_ready),
		.out0(_arith_index_cast3_out0),
		.out0_valid(_arith_index_cast3_out0_valid)
	);
	handshake_buffer_in_ui10_out_ui10_2slots_seq handshake_buffer24(
		.in0(_arith_index_cast3_out0),
		.in0_valid(_arith_index_cast3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(in2_ld0_addr_ready),
		.in0_ready(_handshake_buffer24_in0_ready),
		.out0(in2_ld0_addr),
		.out0_valid(in2_ld0_addr_valid)
	);
	handshake_constant_c0_out_ui64 handshake_constant0(
		.ctrl_valid(_handshake_buffer9_out0_valid),
		.out0_ready(_handshake_buffer25_in0_ready),
		.ctrl_ready(_handshake_constant0_ctrl_ready),
		.out0(_handshake_constant0_out0),
		.out0_valid(_handshake_constant0_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer25(
		.in0(_handshake_constant0_out0),
		.in0_valid(_handshake_constant0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux1_in0_ready),
		.in0_ready(_handshake_buffer25_in0_ready),
		.out0(_handshake_buffer25_out0),
		.out0_valid(_handshake_buffer25_out0_valid)
	);
	handshake_constant_c20_out_ui64 handshake_constant1(
		.ctrl_valid(_handshake_buffer8_out0_valid),
		.out0_ready(_handshake_buffer26_in0_ready),
		.ctrl_ready(_handshake_constant1_ctrl_ready),
		.out0(_handshake_constant1_out0),
		.out0_valid(_handshake_constant1_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer26(
		.in0(_handshake_constant1_out0),
		.in0_valid(_handshake_constant1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux4_in0_ready),
		.in0_ready(_handshake_buffer26_in0_ready),
		.out0(_handshake_buffer26_out0),
		.out0_valid(_handshake_buffer26_out0_valid)
	);
	handshake_constant_c1_out_ui64 handshake_constant2(
		.ctrl_valid(_handshake_buffer7_out0_valid),
		.out0_ready(_handshake_buffer27_in0_ready),
		.ctrl_ready(_handshake_constant2_ctrl_ready),
		.out0(_handshake_constant2_out0),
		.out0_valid(_handshake_constant2_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer27(
		.in0(_handshake_constant2_out0),
		.in0_valid(_handshake_constant2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux5_in0_ready),
		.in0_ready(_handshake_buffer27_in0_ready),
		.out0(_handshake_buffer27_out0),
		.out0_valid(_handshake_buffer27_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_1slots_seq_init_0 handshake_buffer28(
		.in0(_handshake_fork7_out0),
		.in0_valid(_handshake_fork7_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork4_in0_ready),
		.in0_ready(_handshake_buffer28_in0_ready),
		.out0(_handshake_buffer28_out0),
		.out0_valid(_handshake_buffer28_out0_valid)
	);
	handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1 handshake_fork4(
		.in0(_handshake_buffer28_out0),
		.in0_valid(_handshake_buffer28_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer34_in0_ready),
		.out1_ready(_handshake_buffer33_in0_ready),
		.out2_ready(_handshake_buffer32_in0_ready),
		.out3_ready(_handshake_buffer31_in0_ready),
		.out4_ready(_handshake_buffer30_in0_ready),
		.out5_ready(_handshake_buffer29_in0_ready),
		.in0_ready(_handshake_fork4_in0_ready),
		.out0(_handshake_fork4_out0),
		.out0_valid(_handshake_fork4_out0_valid),
		.out1(_handshake_fork4_out1),
		.out1_valid(_handshake_fork4_out1_valid),
		.out2(_handshake_fork4_out2),
		.out2_valid(_handshake_fork4_out2_valid),
		.out3(_handshake_fork4_out3),
		.out3_valid(_handshake_fork4_out3_valid),
		.out4(_handshake_fork4_out4),
		.out4_valid(_handshake_fork4_out4_valid),
		.out5(_handshake_fork4_out5),
		.out5_valid(_handshake_fork4_out5_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer29(
		.in0(_handshake_fork4_out5),
		.in0_valid(_handshake_fork4_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux0_select_ready),
		.in0_ready(_handshake_buffer29_in0_ready),
		.out0(_handshake_buffer29_out0),
		.out0_valid(_handshake_buffer29_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer30(
		.in0(_handshake_fork4_out4),
		.in0_valid(_handshake_fork4_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux1_select_ready),
		.in0_ready(_handshake_buffer30_in0_ready),
		.out0(_handshake_buffer30_out0),
		.out0_valid(_handshake_buffer30_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer31(
		.in0(_handshake_fork4_out3),
		.in0_valid(_handshake_fork4_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux2_select_ready),
		.in0_ready(_handshake_buffer31_in0_ready),
		.out0(_handshake_buffer31_out0),
		.out0_valid(_handshake_buffer31_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer32(
		.in0(_handshake_fork4_out2),
		.in0_valid(_handshake_fork4_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux3_select_ready),
		.in0_ready(_handshake_buffer32_in0_ready),
		.out0(_handshake_buffer32_out0),
		.out0_valid(_handshake_buffer32_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer33(
		.in0(_handshake_fork4_out1),
		.in0_valid(_handshake_fork4_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux4_select_ready),
		.in0_ready(_handshake_buffer33_in0_ready),
		.out0(_handshake_buffer33_out0),
		.out0_valid(_handshake_buffer33_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer34(
		.in0(_handshake_fork4_out0),
		.in0_valid(_handshake_fork4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux5_select_ready),
		.in0_ready(_handshake_buffer34_in0_ready),
		.out0(_handshake_buffer34_out0),
		.out0_valid(_handshake_buffer34_out0_valid)
	);
	handshake_mux_in_ui1_3ins_1outs_ctrl handshake_mux0(
		.select(_handshake_buffer29_out0),
		.select_valid(_handshake_buffer29_out0_valid),
		.in0_valid(_handshake_buffer10_out0_valid),
		.in1_valid(_handshake_buffer119_out0_valid),
		.out0_ready(_handshake_buffer35_in0_ready),
		.select_ready(_handshake_mux0_select_ready),
		.in0_ready(_handshake_mux0_in0_ready),
		.in1_ready(_handshake_mux0_in1_ready),
		.out0_valid(_handshake_mux0_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer35(
		.in0_valid(_handshake_mux0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br5_data_ready),
		.in0_ready(_handshake_buffer35_in0_ready),
		.out0_valid(_handshake_buffer35_out0_valid)
	);
	handshake_mux_in_ui1_ui64_ui64_out_ui64 handshake_mux1(
		.select(_handshake_buffer30_out0),
		.select_valid(_handshake_buffer30_out0_valid),
		.in0(_handshake_buffer25_out0),
		.in0_valid(_handshake_buffer25_out0_valid),
		.in1(_handshake_buffer251_out0),
		.in1_valid(_handshake_buffer251_out0_valid),
		.out0_ready(_handshake_buffer36_in0_ready),
		.select_ready(_handshake_mux1_select_ready),
		.in0_ready(_handshake_mux1_in0_ready),
		.in1_ready(_handshake_mux1_in1_ready),
		.out0(_handshake_mux1_out0),
		.out0_valid(_handshake_mux1_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer36(
		.in0(_handshake_mux1_out0),
		.in0_valid(_handshake_mux1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork5_in0_ready),
		.in0_ready(_handshake_buffer36_in0_ready),
		.out0(_handshake_buffer36_out0),
		.out0_valid(_handshake_buffer36_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork5(
		.in0(_handshake_buffer36_out0),
		.in0_valid(_handshake_buffer36_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer38_in0_ready),
		.out1_ready(_handshake_buffer37_in0_ready),
		.in0_ready(_handshake_fork5_in0_ready),
		.out0(_handshake_fork5_out0),
		.out0_valid(_handshake_fork5_out0_valid),
		.out1(_handshake_fork5_out1),
		.out1_valid(_handshake_fork5_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer37(
		.in0(_handshake_fork5_out1),
		.in0_valid(_handshake_fork5_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br0_data_ready),
		.in0_ready(_handshake_buffer37_in0_ready),
		.out0(_handshake_buffer37_out0),
		.out0_valid(_handshake_buffer37_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer38(
		.in0(_handshake_fork5_out0),
		.in0_valid(_handshake_fork5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi0_in0_ready),
		.in0_ready(_handshake_buffer38_in0_ready),
		.out0(_handshake_buffer38_out0),
		.out0_valid(_handshake_buffer38_out0_valid)
	);
	handshake_mux_in_ui1_ui32_ui32_out_ui32 handshake_mux2(
		.select(_handshake_buffer31_out0),
		.select_valid(_handshake_buffer31_out0_valid),
		.in0(_handshake_buffer6_out0),
		.in0_valid(_handshake_buffer6_out0_valid),
		.in1(_handshake_buffer101_out0),
		.in1_valid(_handshake_buffer101_out0_valid),
		.out0_ready(_handshake_buffer39_in0_ready),
		.select_ready(_handshake_mux2_select_ready),
		.in0_ready(_handshake_mux2_in0_ready),
		.in1_ready(_handshake_mux2_in1_ready),
		.out0(_handshake_mux2_out0),
		.out0_valid(_handshake_mux2_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer39(
		.in0(_handshake_mux2_out0),
		.in0_valid(_handshake_mux2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br1_data_ready),
		.in0_ready(_handshake_buffer39_in0_ready),
		.out0(_handshake_buffer39_out0),
		.out0_valid(_handshake_buffer39_out0_valid)
	);
	handshake_mux_in_ui1_ui32_ui32_out_ui32 handshake_mux3(
		.select(_handshake_buffer32_out0),
		.select_valid(_handshake_buffer32_out0_valid),
		.in0(_handshake_buffer5_out0),
		.in0_valid(_handshake_buffer5_out0_valid),
		.in1(_handshake_buffer103_out0),
		.in1_valid(_handshake_buffer103_out0_valid),
		.out0_ready(_handshake_buffer40_in0_ready),
		.select_ready(_handshake_mux3_select_ready),
		.in0_ready(_handshake_mux3_in0_ready),
		.in1_ready(_handshake_mux3_in1_ready),
		.out0(_handshake_mux3_out0),
		.out0_valid(_handshake_mux3_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer40(
		.in0(_handshake_mux3_out0),
		.in0_valid(_handshake_mux3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br2_data_ready),
		.in0_ready(_handshake_buffer40_in0_ready),
		.out0(_handshake_buffer40_out0),
		.out0_valid(_handshake_buffer40_out0_valid)
	);
	handshake_mux_in_ui1_ui64_ui64_out_ui64 handshake_mux4(
		.select(_handshake_buffer33_out0),
		.select_valid(_handshake_buffer33_out0_valid),
		.in0(_handshake_buffer26_out0),
		.in0_valid(_handshake_buffer26_out0_valid),
		.in1(_handshake_buffer107_out0),
		.in1_valid(_handshake_buffer107_out0_valid),
		.out0_ready(_handshake_buffer41_in0_ready),
		.select_ready(_handshake_mux4_select_ready),
		.in0_ready(_handshake_mux4_in0_ready),
		.in1_ready(_handshake_mux4_in1_ready),
		.out0(_handshake_mux4_out0),
		.out0_valid(_handshake_mux4_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer41(
		.in0(_handshake_mux4_out0),
		.in0_valid(_handshake_mux4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork6_in0_ready),
		.in0_ready(_handshake_buffer41_in0_ready),
		.out0(_handshake_buffer41_out0),
		.out0_valid(_handshake_buffer41_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork6(
		.in0(_handshake_buffer41_out0),
		.in0_valid(_handshake_buffer41_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer43_in0_ready),
		.out1_ready(_handshake_buffer42_in0_ready),
		.in0_ready(_handshake_fork6_in0_ready),
		.out0(_handshake_fork6_out0),
		.out0_valid(_handshake_fork6_out0_valid),
		.out1(_handshake_fork6_out1),
		.out1_valid(_handshake_fork6_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer42(
		.in0(_handshake_fork6_out1),
		.in0_valid(_handshake_fork6_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br3_data_ready),
		.in0_ready(_handshake_buffer42_in0_ready),
		.out0(_handshake_buffer42_out0),
		.out0_valid(_handshake_buffer42_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer43(
		.in0(_handshake_fork6_out0),
		.in0_valid(_handshake_fork6_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi0_in1_ready),
		.in0_ready(_handshake_buffer43_in0_ready),
		.out0(_handshake_buffer43_out0),
		.out0_valid(_handshake_buffer43_out0_valid)
	);
	handshake_mux_in_ui1_ui64_ui64_out_ui64 handshake_mux5(
		.select(_handshake_buffer34_out0),
		.select_valid(_handshake_buffer34_out0_valid),
		.in0(_handshake_buffer27_out0),
		.in0_valid(_handshake_buffer27_out0_valid),
		.in1(_handshake_buffer112_out0),
		.in1_valid(_handshake_buffer112_out0_valid),
		.out0_ready(_handshake_buffer44_in0_ready),
		.select_ready(_handshake_mux5_select_ready),
		.in0_ready(_handshake_mux5_in0_ready),
		.in1_ready(_handshake_mux5_in1_ready),
		.out0(_handshake_mux5_out0),
		.out0_valid(_handshake_mux5_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer44(
		.in0(_handshake_mux5_out0),
		.in0_valid(_handshake_mux5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br4_data_ready),
		.in0_ready(_handshake_buffer44_in0_ready),
		.out0(_handshake_buffer44_out0),
		.out0_valid(_handshake_buffer44_out0_valid)
	);
	arith_cmpi_in_ui64_ui64_out_ui1_slt arith_cmpi0(
		.in0(_handshake_buffer38_out0),
		.in0_valid(_handshake_buffer38_out0_valid),
		.in1(_handshake_buffer43_out0),
		.in1_valid(_handshake_buffer43_out0_valid),
		.out0_ready(_handshake_buffer45_in0_ready),
		.in0_ready(_arith_cmpi0_in0_ready),
		.in1_ready(_arith_cmpi0_in1_ready),
		.out0(_arith_cmpi0_out0),
		.out0_valid(_arith_cmpi0_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer45(
		.in0(_arith_cmpi0_out0),
		.in0_valid(_arith_cmpi0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork7_in0_ready),
		.in0_ready(_handshake_buffer45_in0_ready),
		.out0(_handshake_buffer45_out0),
		.out0_valid(_handshake_buffer45_out0_valid)
	);
	handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1 handshake_fork7(
		.in0(_handshake_buffer45_out0),
		.in0_valid(_handshake_buffer45_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer28_in0_ready),
		.out1_ready(_handshake_buffer51_in0_ready),
		.out2_ready(_handshake_buffer50_in0_ready),
		.out3_ready(_handshake_buffer49_in0_ready),
		.out4_ready(_handshake_buffer48_in0_ready),
		.out5_ready(_handshake_buffer47_in0_ready),
		.out6_ready(_handshake_buffer46_in0_ready),
		.in0_ready(_handshake_fork7_in0_ready),
		.out0(_handshake_fork7_out0),
		.out0_valid(_handshake_fork7_out0_valid),
		.out1(_handshake_fork7_out1),
		.out1_valid(_handshake_fork7_out1_valid),
		.out2(_handshake_fork7_out2),
		.out2_valid(_handshake_fork7_out2_valid),
		.out3(_handshake_fork7_out3),
		.out3_valid(_handshake_fork7_out3_valid),
		.out4(_handshake_fork7_out4),
		.out4_valid(_handshake_fork7_out4_valid),
		.out5(_handshake_fork7_out5),
		.out5_valid(_handshake_fork7_out5_valid),
		.out6(_handshake_fork7_out6),
		.out6_valid(_handshake_fork7_out6_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer46(
		.in0(_handshake_fork7_out6),
		.in0_valid(_handshake_fork7_out6_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br0_cond_ready),
		.in0_ready(_handshake_buffer46_in0_ready),
		.out0(_handshake_buffer46_out0),
		.out0_valid(_handshake_buffer46_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer47(
		.in0(_handshake_fork7_out5),
		.in0_valid(_handshake_fork7_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br1_cond_ready),
		.in0_ready(_handshake_buffer47_in0_ready),
		.out0(_handshake_buffer47_out0),
		.out0_valid(_handshake_buffer47_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer48(
		.in0(_handshake_fork7_out4),
		.in0_valid(_handshake_fork7_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br2_cond_ready),
		.in0_ready(_handshake_buffer48_in0_ready),
		.out0(_handshake_buffer48_out0),
		.out0_valid(_handshake_buffer48_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer49(
		.in0(_handshake_fork7_out3),
		.in0_valid(_handshake_fork7_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br3_cond_ready),
		.in0_ready(_handshake_buffer49_in0_ready),
		.out0(_handshake_buffer49_out0),
		.out0_valid(_handshake_buffer49_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer50(
		.in0(_handshake_fork7_out2),
		.in0_valid(_handshake_fork7_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br4_cond_ready),
		.in0_ready(_handshake_buffer50_in0_ready),
		.out0(_handshake_buffer50_out0),
		.out0_valid(_handshake_buffer50_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer51(
		.in0(_handshake_fork7_out1),
		.in0_valid(_handshake_fork7_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br5_cond_ready),
		.in0_ready(_handshake_buffer51_in0_ready),
		.out0(_handshake_buffer51_out0),
		.out0_valid(_handshake_buffer51_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br0(
		.cond(_handshake_buffer46_out0),
		.cond_valid(_handshake_buffer46_out0_valid),
		.data(_handshake_buffer37_out0),
		.data_valid(_handshake_buffer37_out0_valid),
		.outTrue_ready(_handshake_buffer52_in0_ready),
		.outFalse_ready(_handshake_sink0_in0_ready),
		.cond_ready(_handshake_cond_br0_cond_ready),
		.data_ready(_handshake_cond_br0_data_ready),
		.outTrue(_handshake_cond_br0_outTrue),
		.outTrue_valid(_handshake_cond_br0_outTrue_valid),
		.outFalse(_handshake_cond_br0_outFalse),
		.outFalse_valid(_handshake_cond_br0_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer52(
		.in0(_handshake_cond_br0_outTrue),
		.in0_valid(_handshake_cond_br0_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux11_in0_ready),
		.in0_ready(_handshake_buffer52_in0_ready),
		.out0(_handshake_buffer52_out0),
		.out0_valid(_handshake_buffer52_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink0(
		.in0(_handshake_cond_br0_outFalse),
		.in0_valid(_handshake_cond_br0_outFalse_valid),
		.in0_ready(_handshake_sink0_in0_ready)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br1(
		.cond(_handshake_buffer47_out0),
		.cond_valid(_handshake_buffer47_out0_valid),
		.data(_handshake_buffer39_out0),
		.data_valid(_handshake_buffer39_out0_valid),
		.outTrue_ready(_handshake_buffer53_in0_ready),
		.outFalse_ready(_handshake_sink1_in0_ready),
		.cond_ready(_handshake_cond_br1_cond_ready),
		.data_ready(_handshake_cond_br1_data_ready),
		.outTrue(_handshake_cond_br1_outTrue),
		.outTrue_valid(_handshake_cond_br1_outTrue_valid),
		.outFalse(_handshake_cond_br1_outFalse),
		.outFalse_valid(_handshake_cond_br1_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer53(
		.in0(_handshake_cond_br1_outTrue),
		.in0_valid(_handshake_cond_br1_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux7_in0_ready),
		.in0_ready(_handshake_buffer53_in0_ready),
		.out0(_handshake_buffer53_out0),
		.out0_valid(_handshake_buffer53_out0_valid)
	);
	handshake_sink_in_ui32 handshake_sink1(
		.in0(_handshake_cond_br1_outFalse),
		.in0_valid(_handshake_cond_br1_outFalse_valid),
		.in0_ready(_handshake_sink1_in0_ready)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br2(
		.cond(_handshake_buffer48_out0),
		.cond_valid(_handshake_buffer48_out0_valid),
		.data(_handshake_buffer40_out0),
		.data_valid(_handshake_buffer40_out0_valid),
		.outTrue_ready(_handshake_buffer54_in0_ready),
		.outFalse_ready(_handshake_sink2_in0_ready),
		.cond_ready(_handshake_cond_br2_cond_ready),
		.data_ready(_handshake_cond_br2_data_ready),
		.outTrue(_handshake_cond_br2_outTrue),
		.outTrue_valid(_handshake_cond_br2_outTrue_valid),
		.outFalse(_handshake_cond_br2_outFalse),
		.outFalse_valid(_handshake_cond_br2_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer54(
		.in0(_handshake_cond_br2_outTrue),
		.in0_valid(_handshake_cond_br2_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux8_in0_ready),
		.in0_ready(_handshake_buffer54_in0_ready),
		.out0(_handshake_buffer54_out0),
		.out0_valid(_handshake_buffer54_out0_valid)
	);
	handshake_sink_in_ui32 handshake_sink2(
		.in0(_handshake_cond_br2_outFalse),
		.in0_valid(_handshake_cond_br2_outFalse_valid),
		.in0_ready(_handshake_sink2_in0_ready)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br3(
		.cond(_handshake_buffer49_out0),
		.cond_valid(_handshake_buffer49_out0_valid),
		.data(_handshake_buffer42_out0),
		.data_valid(_handshake_buffer42_out0_valid),
		.outTrue_ready(_handshake_buffer55_in0_ready),
		.outFalse_ready(_handshake_sink3_in0_ready),
		.cond_ready(_handshake_cond_br3_cond_ready),
		.data_ready(_handshake_cond_br3_data_ready),
		.outTrue(_handshake_cond_br3_outTrue),
		.outTrue_valid(_handshake_cond_br3_outTrue_valid),
		.outFalse(_handshake_cond_br3_outFalse),
		.outFalse_valid(_handshake_cond_br3_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer55(
		.in0(_handshake_cond_br3_outTrue),
		.in0_valid(_handshake_cond_br3_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux9_in0_ready),
		.in0_ready(_handshake_buffer55_in0_ready),
		.out0(_handshake_buffer55_out0),
		.out0_valid(_handshake_buffer55_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink3(
		.in0(_handshake_cond_br3_outFalse),
		.in0_valid(_handshake_cond_br3_outFalse_valid),
		.in0_ready(_handshake_sink3_in0_ready)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br4(
		.cond(_handshake_buffer50_out0),
		.cond_valid(_handshake_buffer50_out0_valid),
		.data(_handshake_buffer44_out0),
		.data_valid(_handshake_buffer44_out0_valid),
		.outTrue_ready(_handshake_buffer56_in0_ready),
		.outFalse_ready(_handshake_sink4_in0_ready),
		.cond_ready(_handshake_cond_br4_cond_ready),
		.data_ready(_handshake_cond_br4_data_ready),
		.outTrue(_handshake_cond_br4_outTrue),
		.outTrue_valid(_handshake_cond_br4_outTrue_valid),
		.outFalse(_handshake_cond_br4_outFalse),
		.outFalse_valid(_handshake_cond_br4_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer56(
		.in0(_handshake_cond_br4_outTrue),
		.in0_valid(_handshake_cond_br4_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux10_in0_ready),
		.in0_ready(_handshake_buffer56_in0_ready),
		.out0(_handshake_buffer56_out0),
		.out0_valid(_handshake_buffer56_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink4(
		.in0(_handshake_cond_br4_outFalse),
		.in0_valid(_handshake_cond_br4_outFalse_valid),
		.in0_ready(_handshake_sink4_in0_ready)
	);
	handshake_cond_br_in_ui1_2ins_2outs_ctrl handshake_cond_br5(
		.cond(_handshake_buffer51_out0),
		.cond_valid(_handshake_buffer51_out0_valid),
		.data_valid(_handshake_buffer35_out0_valid),
		.outTrue_ready(_handshake_buffer58_in0_ready),
		.outFalse_ready(_handshake_buffer57_in0_ready),
		.cond_ready(_handshake_cond_br5_cond_ready),
		.data_ready(_handshake_cond_br5_data_ready),
		.outTrue_valid(_handshake_cond_br5_outTrue_valid),
		.outFalse_valid(_handshake_cond_br5_outFalse_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer57(
		.in0_valid(_handshake_cond_br5_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(out0_ready),
		.in0_ready(_handshake_buffer57_in0_ready),
		.out0_valid(out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer58(
		.in0_valid(_handshake_cond_br5_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork8_in0_ready),
		.in0_ready(_handshake_buffer58_in0_ready),
		.out0_valid(_handshake_buffer58_out0_valid)
	);
	handshake_fork_1ins_4outs_ctrl handshake_fork8(
		.in0_valid(_handshake_buffer58_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer62_in0_ready),
		.out1_ready(_handshake_buffer61_in0_ready),
		.out2_ready(_handshake_buffer60_in0_ready),
		.out3_ready(_handshake_buffer59_in0_ready),
		.in0_ready(_handshake_fork8_in0_ready),
		.out0_valid(_handshake_fork8_out0_valid),
		.out1_valid(_handshake_fork8_out1_valid),
		.out2_valid(_handshake_fork8_out2_valid),
		.out3_valid(_handshake_fork8_out3_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer59(
		.in0_valid(_handshake_fork8_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant3_ctrl_ready),
		.in0_ready(_handshake_buffer59_in0_ready),
		.out0_valid(_handshake_buffer59_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer60(
		.in0_valid(_handshake_fork8_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant4_ctrl_ready),
		.in0_ready(_handshake_buffer60_in0_ready),
		.out0_valid(_handshake_buffer60_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer61(
		.in0_valid(_handshake_fork8_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant5_ctrl_ready),
		.in0_ready(_handshake_buffer61_in0_ready),
		.out0_valid(_handshake_buffer61_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer62(
		.in0_valid(_handshake_fork8_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_control_merge0_in0_ready),
		.in0_ready(_handshake_buffer62_in0_ready),
		.out0_valid(_handshake_buffer62_out0_valid)
	);
	handshake_constant_c0_out_ui64 handshake_constant3(
		.ctrl_valid(_handshake_buffer59_out0_valid),
		.out0_ready(_handshake_buffer63_in0_ready),
		.ctrl_ready(_handshake_constant3_ctrl_ready),
		.out0(_handshake_constant3_out0),
		.out0_valid(_handshake_constant3_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer63(
		.in0(_handshake_constant3_out0),
		.in0_valid(_handshake_constant3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux6_in0_ready),
		.in0_ready(_handshake_buffer63_in0_ready),
		.out0(_handshake_buffer63_out0),
		.out0_valid(_handshake_buffer63_out0_valid)
	);
	handshake_constant_c20_out_ui64 handshake_constant4(
		.ctrl_valid(_handshake_buffer60_out0_valid),
		.out0_ready(_handshake_buffer64_in0_ready),
		.ctrl_ready(_handshake_constant4_ctrl_ready),
		.out0(_handshake_constant4_out0),
		.out0_valid(_handshake_constant4_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer64(
		.in0(_handshake_constant4_out0),
		.in0_valid(_handshake_constant4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux12_in0_ready),
		.in0_ready(_handshake_buffer64_in0_ready),
		.out0(_handshake_buffer64_out0),
		.out0_valid(_handshake_buffer64_out0_valid)
	);
	handshake_constant_c1_out_ui64 handshake_constant5(
		.ctrl_valid(_handshake_buffer61_out0_valid),
		.out0_ready(_handshake_buffer65_in0_ready),
		.ctrl_ready(_handshake_constant5_ctrl_ready),
		.out0(_handshake_constant5_out0),
		.out0_valid(_handshake_constant5_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer65(
		.in0(_handshake_constant5_out0),
		.in0_valid(_handshake_constant5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux13_in0_ready),
		.in0_ready(_handshake_buffer65_in0_ready),
		.out0(_handshake_buffer65_out0),
		.out0_valid(_handshake_buffer65_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux6(
		.select(_handshake_buffer80_out0),
		.select_valid(_handshake_buffer80_out0_valid),
		.in0(_handshake_buffer63_out0),
		.in0_valid(_handshake_buffer63_out0_valid),
		.in1(_handshake_buffer250_out0),
		.in1_valid(_handshake_buffer250_out0_valid),
		.out0_ready(_handshake_buffer66_in0_ready),
		.select_ready(_handshake_mux6_select_ready),
		.in0_ready(_handshake_mux6_in0_ready),
		.in1_ready(_handshake_mux6_in1_ready),
		.out0(_handshake_mux6_out0),
		.out0_valid(_handshake_mux6_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer66(
		.in0(_handshake_mux6_out0),
		.in0_valid(_handshake_mux6_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork9_in0_ready),
		.in0_ready(_handshake_buffer66_in0_ready),
		.out0(_handshake_buffer66_out0),
		.out0_valid(_handshake_buffer66_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork9(
		.in0(_handshake_buffer66_out0),
		.in0_valid(_handshake_buffer66_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer68_in0_ready),
		.out1_ready(_handshake_buffer67_in0_ready),
		.in0_ready(_handshake_fork9_in0_ready),
		.out0(_handshake_fork9_out0),
		.out0_valid(_handshake_fork9_out0_valid),
		.out1(_handshake_fork9_out1),
		.out1_valid(_handshake_fork9_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer67(
		.in0(_handshake_fork9_out1),
		.in0_valid(_handshake_fork9_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi1_in0_ready),
		.in0_ready(_handshake_buffer67_in0_ready),
		.out0(_handshake_buffer67_out0),
		.out0_valid(_handshake_buffer67_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer68(
		.in0(_handshake_fork9_out0),
		.in0_valid(_handshake_fork9_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br6_data_ready),
		.in0_ready(_handshake_buffer68_in0_ready),
		.out0(_handshake_buffer68_out0),
		.out0_valid(_handshake_buffer68_out0_valid)
	);
	handshake_mux_in_ui64_ui32_ui32_out_ui32 handshake_mux7(
		.select(_handshake_buffer81_out0),
		.select_valid(_handshake_buffer81_out0_valid),
		.in0(_handshake_buffer53_out0),
		.in0_valid(_handshake_buffer53_out0_valid),
		.in1(_handshake_buffer187_out0),
		.in1_valid(_handshake_buffer187_out0_valid),
		.out0_ready(_handshake_buffer69_in0_ready),
		.select_ready(_handshake_mux7_select_ready),
		.in0_ready(_handshake_mux7_in0_ready),
		.in1_ready(_handshake_mux7_in1_ready),
		.out0(_handshake_mux7_out0),
		.out0_valid(_handshake_mux7_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer69(
		.in0(_handshake_mux7_out0),
		.in0_valid(_handshake_mux7_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br7_data_ready),
		.in0_ready(_handshake_buffer69_in0_ready),
		.out0(_handshake_buffer69_out0),
		.out0_valid(_handshake_buffer69_out0_valid)
	);
	handshake_mux_in_ui64_ui32_ui32_out_ui32 handshake_mux8(
		.select(_handshake_buffer82_out0),
		.select_valid(_handshake_buffer82_out0_valid),
		.in0(_handshake_buffer54_out0),
		.in0_valid(_handshake_buffer54_out0_valid),
		.in1(_handshake_buffer191_out0),
		.in1_valid(_handshake_buffer191_out0_valid),
		.out0_ready(_handshake_buffer70_in0_ready),
		.select_ready(_handshake_mux8_select_ready),
		.in0_ready(_handshake_mux8_in0_ready),
		.in1_ready(_handshake_mux8_in1_ready),
		.out0(_handshake_mux8_out0),
		.out0_valid(_handshake_mux8_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer70(
		.in0(_handshake_mux8_out0),
		.in0_valid(_handshake_mux8_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br8_data_ready),
		.in0_ready(_handshake_buffer70_in0_ready),
		.out0(_handshake_buffer70_out0),
		.out0_valid(_handshake_buffer70_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux9(
		.select(_handshake_buffer83_out0),
		.select_valid(_handshake_buffer83_out0_valid),
		.in0(_handshake_buffer55_out0),
		.in0_valid(_handshake_buffer55_out0_valid),
		.in1(_handshake_buffer193_out0),
		.in1_valid(_handshake_buffer193_out0_valid),
		.out0_ready(_handshake_buffer71_in0_ready),
		.select_ready(_handshake_mux9_select_ready),
		.in0_ready(_handshake_mux9_in0_ready),
		.in1_ready(_handshake_mux9_in1_ready),
		.out0(_handshake_mux9_out0),
		.out0_valid(_handshake_mux9_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer71(
		.in0(_handshake_mux9_out0),
		.in0_valid(_handshake_mux9_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br9_data_ready),
		.in0_ready(_handshake_buffer71_in0_ready),
		.out0(_handshake_buffer71_out0),
		.out0_valid(_handshake_buffer71_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux10(
		.select(_handshake_buffer84_out0),
		.select_valid(_handshake_buffer84_out0_valid),
		.in0(_handshake_buffer56_out0),
		.in0_valid(_handshake_buffer56_out0_valid),
		.in1(_handshake_buffer195_out0),
		.in1_valid(_handshake_buffer195_out0_valid),
		.out0_ready(_handshake_buffer72_in0_ready),
		.select_ready(_handshake_mux10_select_ready),
		.in0_ready(_handshake_mux10_in0_ready),
		.in1_ready(_handshake_mux10_in1_ready),
		.out0(_handshake_mux10_out0),
		.out0_valid(_handshake_mux10_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer72(
		.in0(_handshake_mux10_out0),
		.in0_valid(_handshake_mux10_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br10_data_ready),
		.in0_ready(_handshake_buffer72_in0_ready),
		.out0(_handshake_buffer72_out0),
		.out0_valid(_handshake_buffer72_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux11(
		.select(_handshake_buffer85_out0),
		.select_valid(_handshake_buffer85_out0_valid),
		.in0(_handshake_buffer52_out0),
		.in0_valid(_handshake_buffer52_out0_valid),
		.in1(_handshake_buffer200_out0),
		.in1_valid(_handshake_buffer200_out0_valid),
		.out0_ready(_handshake_buffer73_in0_ready),
		.select_ready(_handshake_mux11_select_ready),
		.in0_ready(_handshake_mux11_in0_ready),
		.in1_ready(_handshake_mux11_in1_ready),
		.out0(_handshake_mux11_out0),
		.out0_valid(_handshake_mux11_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer73(
		.in0(_handshake_mux11_out0),
		.in0_valid(_handshake_mux11_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br11_data_ready),
		.in0_ready(_handshake_buffer73_in0_ready),
		.out0(_handshake_buffer73_out0),
		.out0_valid(_handshake_buffer73_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux12(
		.select(_handshake_buffer86_out0),
		.select_valid(_handshake_buffer86_out0_valid),
		.in0(_handshake_buffer64_out0),
		.in0_valid(_handshake_buffer64_out0_valid),
		.in1(_handshake_buffer203_out0),
		.in1_valid(_handshake_buffer203_out0_valid),
		.out0_ready(_handshake_buffer74_in0_ready),
		.select_ready(_handshake_mux12_select_ready),
		.in0_ready(_handshake_mux12_in0_ready),
		.in1_ready(_handshake_mux12_in1_ready),
		.out0(_handshake_mux12_out0),
		.out0_valid(_handshake_mux12_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer74(
		.in0(_handshake_mux12_out0),
		.in0_valid(_handshake_mux12_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork10_in0_ready),
		.in0_ready(_handshake_buffer74_in0_ready),
		.out0(_handshake_buffer74_out0),
		.out0_valid(_handshake_buffer74_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork10(
		.in0(_handshake_buffer74_out0),
		.in0_valid(_handshake_buffer74_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer76_in0_ready),
		.out1_ready(_handshake_buffer75_in0_ready),
		.in0_ready(_handshake_fork10_in0_ready),
		.out0(_handshake_fork10_out0),
		.out0_valid(_handshake_fork10_out0_valid),
		.out1(_handshake_fork10_out1),
		.out1_valid(_handshake_fork10_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer75(
		.in0(_handshake_fork10_out1),
		.in0_valid(_handshake_fork10_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi1_in1_ready),
		.in0_ready(_handshake_buffer75_in0_ready),
		.out0(_handshake_buffer75_out0),
		.out0_valid(_handshake_buffer75_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer76(
		.in0(_handshake_fork10_out0),
		.in0_valid(_handshake_fork10_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br12_data_ready),
		.in0_ready(_handshake_buffer76_in0_ready),
		.out0(_handshake_buffer76_out0),
		.out0_valid(_handshake_buffer76_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux13(
		.select(_handshake_buffer87_out0),
		.select_valid(_handshake_buffer87_out0_valid),
		.in0(_handshake_buffer65_out0),
		.in0_valid(_handshake_buffer65_out0_valid),
		.in1(_handshake_buffer208_out0),
		.in1_valid(_handshake_buffer208_out0_valid),
		.out0_ready(_handshake_buffer77_in0_ready),
		.select_ready(_handshake_mux13_select_ready),
		.in0_ready(_handshake_mux13_in0_ready),
		.in1_ready(_handshake_mux13_in1_ready),
		.out0(_handshake_mux13_out0),
		.out0_valid(_handshake_mux13_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer77(
		.in0(_handshake_mux13_out0),
		.in0_valid(_handshake_mux13_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br13_data_ready),
		.in0_ready(_handshake_buffer77_in0_ready),
		.out0(_handshake_buffer77_out0),
		.out0_valid(_handshake_buffer77_out0_valid)
	);
	handshake_control_merge_out_ui64_2ins_2outs_ctrl handshake_control_merge0(
		.in0_valid(_handshake_buffer62_out0_valid),
		.in1_valid(_handshake_buffer244_out0_valid),
		.clock(clock),
		.reset(reset),
		.dataOut_ready(_handshake_buffer79_in0_ready),
		.index_ready(_handshake_buffer78_in0_ready),
		.in0_ready(_handshake_control_merge0_in0_ready),
		.in1_ready(_handshake_control_merge0_in1_ready),
		.dataOut_valid(_handshake_control_merge0_dataOut_valid),
		.index(_handshake_control_merge0_index),
		.index_valid(_handshake_control_merge0_index_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer78(
		.in0(_handshake_control_merge0_index),
		.in0_valid(_handshake_control_merge0_index_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork11_in0_ready),
		.in0_ready(_handshake_buffer78_in0_ready),
		.out0(_handshake_buffer78_out0),
		.out0_valid(_handshake_buffer78_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer79(
		.in0_valid(_handshake_control_merge0_dataOut_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br14_data_ready),
		.in0_ready(_handshake_buffer79_in0_ready),
		.out0_valid(_handshake_buffer79_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64 handshake_fork11(
		.in0(_handshake_buffer78_out0),
		.in0_valid(_handshake_buffer78_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer87_in0_ready),
		.out1_ready(_handshake_buffer86_in0_ready),
		.out2_ready(_handshake_buffer85_in0_ready),
		.out3_ready(_handshake_buffer84_in0_ready),
		.out4_ready(_handshake_buffer83_in0_ready),
		.out5_ready(_handshake_buffer82_in0_ready),
		.out6_ready(_handshake_buffer81_in0_ready),
		.out7_ready(_handshake_buffer80_in0_ready),
		.in0_ready(_handshake_fork11_in0_ready),
		.out0(_handshake_fork11_out0),
		.out0_valid(_handshake_fork11_out0_valid),
		.out1(_handshake_fork11_out1),
		.out1_valid(_handshake_fork11_out1_valid),
		.out2(_handshake_fork11_out2),
		.out2_valid(_handshake_fork11_out2_valid),
		.out3(_handshake_fork11_out3),
		.out3_valid(_handshake_fork11_out3_valid),
		.out4(_handshake_fork11_out4),
		.out4_valid(_handshake_fork11_out4_valid),
		.out5(_handshake_fork11_out5),
		.out5_valid(_handshake_fork11_out5_valid),
		.out6(_handshake_fork11_out6),
		.out6_valid(_handshake_fork11_out6_valid),
		.out7(_handshake_fork11_out7),
		.out7_valid(_handshake_fork11_out7_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer80(
		.in0(_handshake_fork11_out7),
		.in0_valid(_handshake_fork11_out7_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux6_select_ready),
		.in0_ready(_handshake_buffer80_in0_ready),
		.out0(_handshake_buffer80_out0),
		.out0_valid(_handshake_buffer80_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer81(
		.in0(_handshake_fork11_out6),
		.in0_valid(_handshake_fork11_out6_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux7_select_ready),
		.in0_ready(_handshake_buffer81_in0_ready),
		.out0(_handshake_buffer81_out0),
		.out0_valid(_handshake_buffer81_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer82(
		.in0(_handshake_fork11_out5),
		.in0_valid(_handshake_fork11_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux8_select_ready),
		.in0_ready(_handshake_buffer82_in0_ready),
		.out0(_handshake_buffer82_out0),
		.out0_valid(_handshake_buffer82_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer83(
		.in0(_handshake_fork11_out4),
		.in0_valid(_handshake_fork11_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux9_select_ready),
		.in0_ready(_handshake_buffer83_in0_ready),
		.out0(_handshake_buffer83_out0),
		.out0_valid(_handshake_buffer83_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer84(
		.in0(_handshake_fork11_out3),
		.in0_valid(_handshake_fork11_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux10_select_ready),
		.in0_ready(_handshake_buffer84_in0_ready),
		.out0(_handshake_buffer84_out0),
		.out0_valid(_handshake_buffer84_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer85(
		.in0(_handshake_fork11_out2),
		.in0_valid(_handshake_fork11_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux11_select_ready),
		.in0_ready(_handshake_buffer85_in0_ready),
		.out0(_handshake_buffer85_out0),
		.out0_valid(_handshake_buffer85_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer86(
		.in0(_handshake_fork11_out1),
		.in0_valid(_handshake_fork11_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux12_select_ready),
		.in0_ready(_handshake_buffer86_in0_ready),
		.out0(_handshake_buffer86_out0),
		.out0_valid(_handshake_buffer86_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer87(
		.in0(_handshake_fork11_out0),
		.in0_valid(_handshake_fork11_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux13_select_ready),
		.in0_ready(_handshake_buffer87_in0_ready),
		.out0(_handshake_buffer87_out0),
		.out0_valid(_handshake_buffer87_out0_valid)
	);
	arith_cmpi_in_ui64_ui64_out_ui1_slt arith_cmpi1(
		.in0(_handshake_buffer67_out0),
		.in0_valid(_handshake_buffer67_out0_valid),
		.in1(_handshake_buffer75_out0),
		.in1_valid(_handshake_buffer75_out0_valid),
		.out0_ready(_handshake_buffer88_in0_ready),
		.in0_ready(_arith_cmpi1_in0_ready),
		.in1_ready(_arith_cmpi1_in1_ready),
		.out0(_arith_cmpi1_out0),
		.out0_valid(_arith_cmpi1_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer88(
		.in0(_arith_cmpi1_out0),
		.in0_valid(_arith_cmpi1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork12_in0_ready),
		.in0_ready(_handshake_buffer88_in0_ready),
		.out0(_handshake_buffer88_out0),
		.out0_valid(_handshake_buffer88_out0_valid)
	);
	handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1 handshake_fork12(
		.in0(_handshake_buffer88_out0),
		.in0_valid(_handshake_buffer88_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer97_in0_ready),
		.out1_ready(_handshake_buffer96_in0_ready),
		.out2_ready(_handshake_buffer95_in0_ready),
		.out3_ready(_handshake_buffer94_in0_ready),
		.out4_ready(_handshake_buffer93_in0_ready),
		.out5_ready(_handshake_buffer92_in0_ready),
		.out6_ready(_handshake_buffer91_in0_ready),
		.out7_ready(_handshake_buffer90_in0_ready),
		.out8_ready(_handshake_buffer89_in0_ready),
		.in0_ready(_handshake_fork12_in0_ready),
		.out0(_handshake_fork12_out0),
		.out0_valid(_handshake_fork12_out0_valid),
		.out1(_handshake_fork12_out1),
		.out1_valid(_handshake_fork12_out1_valid),
		.out2(_handshake_fork12_out2),
		.out2_valid(_handshake_fork12_out2_valid),
		.out3(_handshake_fork12_out3),
		.out3_valid(_handshake_fork12_out3_valid),
		.out4(_handshake_fork12_out4),
		.out4_valid(_handshake_fork12_out4_valid),
		.out5(_handshake_fork12_out5),
		.out5_valid(_handshake_fork12_out5_valid),
		.out6(_handshake_fork12_out6),
		.out6_valid(_handshake_fork12_out6_valid),
		.out7(_handshake_fork12_out7),
		.out7_valid(_handshake_fork12_out7_valid),
		.out8(_handshake_fork12_out8),
		.out8_valid(_handshake_fork12_out8_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer89(
		.in0(_handshake_fork12_out8),
		.in0_valid(_handshake_fork12_out8_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br6_cond_ready),
		.in0_ready(_handshake_buffer89_in0_ready),
		.out0(_handshake_buffer89_out0),
		.out0_valid(_handshake_buffer89_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer90(
		.in0(_handshake_fork12_out7),
		.in0_valid(_handshake_fork12_out7_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br7_cond_ready),
		.in0_ready(_handshake_buffer90_in0_ready),
		.out0(_handshake_buffer90_out0),
		.out0_valid(_handshake_buffer90_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer91(
		.in0(_handshake_fork12_out6),
		.in0_valid(_handshake_fork12_out6_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br8_cond_ready),
		.in0_ready(_handshake_buffer91_in0_ready),
		.out0(_handshake_buffer91_out0),
		.out0_valid(_handshake_buffer91_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer92(
		.in0(_handshake_fork12_out5),
		.in0_valid(_handshake_fork12_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br9_cond_ready),
		.in0_ready(_handshake_buffer92_in0_ready),
		.out0(_handshake_buffer92_out0),
		.out0_valid(_handshake_buffer92_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer93(
		.in0(_handshake_fork12_out4),
		.in0_valid(_handshake_fork12_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br10_cond_ready),
		.in0_ready(_handshake_buffer93_in0_ready),
		.out0(_handshake_buffer93_out0),
		.out0_valid(_handshake_buffer93_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer94(
		.in0(_handshake_fork12_out3),
		.in0_valid(_handshake_fork12_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br11_cond_ready),
		.in0_ready(_handshake_buffer94_in0_ready),
		.out0(_handshake_buffer94_out0),
		.out0_valid(_handshake_buffer94_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer95(
		.in0(_handshake_fork12_out2),
		.in0_valid(_handshake_fork12_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br12_cond_ready),
		.in0_ready(_handshake_buffer95_in0_ready),
		.out0(_handshake_buffer95_out0),
		.out0_valid(_handshake_buffer95_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer96(
		.in0(_handshake_fork12_out1),
		.in0_valid(_handshake_fork12_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br13_cond_ready),
		.in0_ready(_handshake_buffer96_in0_ready),
		.out0(_handshake_buffer96_out0),
		.out0_valid(_handshake_buffer96_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer97(
		.in0(_handshake_fork12_out0),
		.in0_valid(_handshake_fork12_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br14_cond_ready),
		.in0_ready(_handshake_buffer97_in0_ready),
		.out0(_handshake_buffer97_out0),
		.out0_valid(_handshake_buffer97_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br6(
		.cond(_handshake_buffer89_out0),
		.cond_valid(_handshake_buffer89_out0_valid),
		.data(_handshake_buffer68_out0),
		.data_valid(_handshake_buffer68_out0_valid),
		.outTrue_ready(_handshake_buffer98_in0_ready),
		.outFalse_ready(_handshake_sink5_in0_ready),
		.cond_ready(_handshake_cond_br6_cond_ready),
		.data_ready(_handshake_cond_br6_data_ready),
		.outTrue(_handshake_cond_br6_outTrue),
		.outTrue_valid(_handshake_cond_br6_outTrue_valid),
		.outFalse(_handshake_cond_br6_outFalse),
		.outFalse_valid(_handshake_cond_br6_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer98(
		.in0(_handshake_cond_br6_outTrue),
		.in0_valid(_handshake_cond_br6_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork13_in0_ready),
		.in0_ready(_handshake_buffer98_in0_ready),
		.out0(_handshake_buffer98_out0),
		.out0_valid(_handshake_buffer98_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink5(
		.in0(_handshake_cond_br6_outFalse),
		.in0_valid(_handshake_cond_br6_outFalse_valid),
		.in0_ready(_handshake_sink5_in0_ready)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork13(
		.in0(_handshake_buffer98_out0),
		.in0_valid(_handshake_buffer98_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer100_in0_ready),
		.out1_ready(_handshake_buffer99_in0_ready),
		.in0_ready(_handshake_fork13_in0_ready),
		.out0(_handshake_fork13_out0),
		.out0_valid(_handshake_fork13_out0_valid),
		.out1(_handshake_fork13_out1),
		.out1_valid(_handshake_fork13_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer99(
		.in0(_handshake_fork13_out1),
		.in0_valid(_handshake_fork13_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi0_in1_ready),
		.in0_ready(_handshake_buffer99_in0_ready),
		.out0(_handshake_buffer99_out0),
		.out0_valid(_handshake_buffer99_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer100(
		.in0(_handshake_fork13_out0),
		.in0_valid(_handshake_fork13_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux23_in0_ready),
		.in0_ready(_handshake_buffer100_in0_ready),
		.out0(_handshake_buffer100_out0),
		.out0_valid(_handshake_buffer100_out0_valid)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br7(
		.cond(_handshake_buffer90_out0),
		.cond_valid(_handshake_buffer90_out0_valid),
		.data(_handshake_buffer69_out0),
		.data_valid(_handshake_buffer69_out0_valid),
		.outTrue_ready(_handshake_buffer102_in0_ready),
		.outFalse_ready(_handshake_buffer101_in0_ready),
		.cond_ready(_handshake_cond_br7_cond_ready),
		.data_ready(_handshake_cond_br7_data_ready),
		.outTrue(_handshake_cond_br7_outTrue),
		.outTrue_valid(_handshake_cond_br7_outTrue_valid),
		.outFalse(_handshake_cond_br7_outFalse),
		.outFalse_valid(_handshake_cond_br7_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer101(
		.in0(_handshake_cond_br7_outFalse),
		.in0_valid(_handshake_cond_br7_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux2_in1_ready),
		.in0_ready(_handshake_buffer101_in0_ready),
		.out0(_handshake_buffer101_out0),
		.out0_valid(_handshake_buffer101_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer102(
		.in0(_handshake_cond_br7_outTrue),
		.in0_valid(_handshake_cond_br7_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux16_in0_ready),
		.in0_ready(_handshake_buffer102_in0_ready),
		.out0(_handshake_buffer102_out0),
		.out0_valid(_handshake_buffer102_out0_valid)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br8(
		.cond(_handshake_buffer91_out0),
		.cond_valid(_handshake_buffer91_out0_valid),
		.data(_handshake_buffer70_out0),
		.data_valid(_handshake_buffer70_out0_valid),
		.outTrue_ready(_handshake_buffer104_in0_ready),
		.outFalse_ready(_handshake_buffer103_in0_ready),
		.cond_ready(_handshake_cond_br8_cond_ready),
		.data_ready(_handshake_cond_br8_data_ready),
		.outTrue(_handshake_cond_br8_outTrue),
		.outTrue_valid(_handshake_cond_br8_outTrue_valid),
		.outFalse(_handshake_cond_br8_outFalse),
		.outFalse_valid(_handshake_cond_br8_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer103(
		.in0(_handshake_cond_br8_outFalse),
		.in0_valid(_handshake_cond_br8_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux3_in1_ready),
		.in0_ready(_handshake_buffer103_in0_ready),
		.out0(_handshake_buffer103_out0),
		.out0_valid(_handshake_buffer103_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer104(
		.in0(_handshake_cond_br8_outTrue),
		.in0_valid(_handshake_cond_br8_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork14_in0_ready),
		.in0_ready(_handshake_buffer104_in0_ready),
		.out0(_handshake_buffer104_out0),
		.out0_valid(_handshake_buffer104_out0_valid)
	);
	handshake_fork_in_ui32_out_ui32_ui32 handshake_fork14(
		.in0(_handshake_buffer104_out0),
		.in0_valid(_handshake_buffer104_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer106_in0_ready),
		.out1_ready(_handshake_buffer105_in0_ready),
		.in0_ready(_handshake_fork14_in0_ready),
		.out0(_handshake_fork14_out0),
		.out0_valid(_handshake_fork14_out0_valid),
		.out1(_handshake_fork14_out1),
		.out1_valid(_handshake_fork14_out1_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer105(
		.in0(_handshake_fork14_out1),
		.in0_valid(_handshake_fork14_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli1_in1_ready),
		.in0_ready(_handshake_buffer105_in0_ready),
		.out0(_handshake_buffer105_out0),
		.out0_valid(_handshake_buffer105_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer106(
		.in0(_handshake_fork14_out0),
		.in0_valid(_handshake_fork14_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux17_in0_ready),
		.in0_ready(_handshake_buffer106_in0_ready),
		.out0(_handshake_buffer106_out0),
		.out0_valid(_handshake_buffer106_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br9(
		.cond(_handshake_buffer92_out0),
		.cond_valid(_handshake_buffer92_out0_valid),
		.data(_handshake_buffer71_out0),
		.data_valid(_handshake_buffer71_out0_valid),
		.outTrue_ready(_handshake_buffer108_in0_ready),
		.outFalse_ready(_handshake_buffer107_in0_ready),
		.cond_ready(_handshake_cond_br9_cond_ready),
		.data_ready(_handshake_cond_br9_data_ready),
		.outTrue(_handshake_cond_br9_outTrue),
		.outTrue_valid(_handshake_cond_br9_outTrue_valid),
		.outFalse(_handshake_cond_br9_outFalse),
		.outFalse_valid(_handshake_cond_br9_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer107(
		.in0(_handshake_cond_br9_outFalse),
		.in0_valid(_handshake_cond_br9_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux4_in1_ready),
		.in0_ready(_handshake_buffer107_in0_ready),
		.out0(_handshake_buffer107_out0),
		.out0_valid(_handshake_buffer107_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer108(
		.in0(_handshake_cond_br9_outTrue),
		.in0_valid(_handshake_cond_br9_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux18_in0_ready),
		.in0_ready(_handshake_buffer108_in0_ready),
		.out0(_handshake_buffer108_out0),
		.out0_valid(_handshake_buffer108_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br10(
		.cond(_handshake_buffer93_out0),
		.cond_valid(_handshake_buffer93_out0_valid),
		.data(_handshake_buffer72_out0),
		.data_valid(_handshake_buffer72_out0_valid),
		.outTrue_ready(_handshake_buffer110_in0_ready),
		.outFalse_ready(_handshake_buffer109_in0_ready),
		.cond_ready(_handshake_cond_br10_cond_ready),
		.data_ready(_handshake_cond_br10_data_ready),
		.outTrue(_handshake_cond_br10_outTrue),
		.outTrue_valid(_handshake_cond_br10_outTrue_valid),
		.outFalse(_handshake_cond_br10_outFalse),
		.outFalse_valid(_handshake_cond_br10_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer109(
		.in0(_handshake_cond_br10_outFalse),
		.in0_valid(_handshake_cond_br10_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork15_in0_ready),
		.in0_ready(_handshake_buffer109_in0_ready),
		.out0(_handshake_buffer109_out0),
		.out0_valid(_handshake_buffer109_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer110(
		.in0(_handshake_cond_br10_outTrue),
		.in0_valid(_handshake_cond_br10_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux19_in0_ready),
		.in0_ready(_handshake_buffer110_in0_ready),
		.out0(_handshake_buffer110_out0),
		.out0_valid(_handshake_buffer110_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork15(
		.in0(_handshake_buffer109_out0),
		.in0_valid(_handshake_buffer109_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer112_in0_ready),
		.out1_ready(_handshake_buffer111_in0_ready),
		.in0_ready(_handshake_fork15_in0_ready),
		.out0(_handshake_fork15_out0),
		.out0_valid(_handshake_fork15_out0_valid),
		.out1(_handshake_fork15_out1),
		.out1_valid(_handshake_fork15_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer111(
		.in0(_handshake_fork15_out1),
		.in0_valid(_handshake_fork15_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi7_in1_ready),
		.in0_ready(_handshake_buffer111_in0_ready),
		.out0(_handshake_buffer111_out0),
		.out0_valid(_handshake_buffer111_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer112(
		.in0(_handshake_fork15_out0),
		.in0_valid(_handshake_fork15_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux5_in1_ready),
		.in0_ready(_handshake_buffer112_in0_ready),
		.out0(_handshake_buffer112_out0),
		.out0_valid(_handshake_buffer112_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br11(
		.cond(_handshake_buffer94_out0),
		.cond_valid(_handshake_buffer94_out0_valid),
		.data(_handshake_buffer73_out0),
		.data_valid(_handshake_buffer73_out0_valid),
		.outTrue_ready(_handshake_buffer114_in0_ready),
		.outFalse_ready(_handshake_buffer113_in0_ready),
		.cond_ready(_handshake_cond_br11_cond_ready),
		.data_ready(_handshake_cond_br11_data_ready),
		.outTrue(_handshake_cond_br11_outTrue),
		.outTrue_valid(_handshake_cond_br11_outTrue_valid),
		.outFalse(_handshake_cond_br11_outFalse),
		.outFalse_valid(_handshake_cond_br11_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer113(
		.in0(_handshake_cond_br11_outFalse),
		.in0_valid(_handshake_cond_br11_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi7_in0_ready),
		.in0_ready(_handshake_buffer113_in0_ready),
		.out0(_handshake_buffer113_out0),
		.out0_valid(_handshake_buffer113_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer114(
		.in0(_handshake_cond_br11_outTrue),
		.in0_valid(_handshake_cond_br11_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork16_in0_ready),
		.in0_ready(_handshake_buffer114_in0_ready),
		.out0(_handshake_buffer114_out0),
		.out0_valid(_handshake_buffer114_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork16(
		.in0(_handshake_buffer114_out0),
		.in0_valid(_handshake_buffer114_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer116_in0_ready),
		.out1_ready(_handshake_buffer115_in0_ready),
		.in0_ready(_handshake_fork16_in0_ready),
		.out0(_handshake_fork16_out0),
		.out0_valid(_handshake_fork16_out0_valid),
		.out1(_handshake_fork16_out1),
		.out1_valid(_handshake_fork16_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer115(
		.in0(_handshake_fork16_out1),
		.in0_valid(_handshake_fork16_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli0_in0_ready),
		.in0_ready(_handshake_buffer115_in0_ready),
		.out0(_handshake_buffer115_out0),
		.out0_valid(_handshake_buffer115_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer116(
		.in0(_handshake_fork16_out0),
		.in0_valid(_handshake_fork16_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux20_in0_ready),
		.in0_ready(_handshake_buffer116_in0_ready),
		.out0(_handshake_buffer116_out0),
		.out0_valid(_handshake_buffer116_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br12(
		.cond(_handshake_buffer95_out0),
		.cond_valid(_handshake_buffer95_out0_valid),
		.data(_handshake_buffer76_out0),
		.data_valid(_handshake_buffer76_out0_valid),
		.outTrue_ready(_handshake_buffer117_in0_ready),
		.outFalse_ready(_handshake_sink6_in0_ready),
		.cond_ready(_handshake_cond_br12_cond_ready),
		.data_ready(_handshake_cond_br12_data_ready),
		.outTrue(_handshake_cond_br12_outTrue),
		.outTrue_valid(_handshake_cond_br12_outTrue_valid),
		.outFalse(_handshake_cond_br12_outFalse),
		.outFalse_valid(_handshake_cond_br12_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer117(
		.in0(_handshake_cond_br12_outTrue),
		.in0_valid(_handshake_cond_br12_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux21_in0_ready),
		.in0_ready(_handshake_buffer117_in0_ready),
		.out0(_handshake_buffer117_out0),
		.out0_valid(_handshake_buffer117_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink6(
		.in0(_handshake_cond_br12_outFalse),
		.in0_valid(_handshake_cond_br12_outFalse_valid),
		.in0_ready(_handshake_sink6_in0_ready)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br13(
		.cond(_handshake_buffer96_out0),
		.cond_valid(_handshake_buffer96_out0_valid),
		.data(_handshake_buffer77_out0),
		.data_valid(_handshake_buffer77_out0_valid),
		.outTrue_ready(_handshake_buffer118_in0_ready),
		.outFalse_ready(_handshake_sink7_in0_ready),
		.cond_ready(_handshake_cond_br13_cond_ready),
		.data_ready(_handshake_cond_br13_data_ready),
		.outTrue(_handshake_cond_br13_outTrue),
		.outTrue_valid(_handshake_cond_br13_outTrue_valid),
		.outFalse(_handshake_cond_br13_outFalse),
		.outFalse_valid(_handshake_cond_br13_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer118(
		.in0(_handshake_cond_br13_outTrue),
		.in0_valid(_handshake_cond_br13_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux22_in0_ready),
		.in0_ready(_handshake_buffer118_in0_ready),
		.out0(_handshake_buffer118_out0),
		.out0_valid(_handshake_buffer118_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink7(
		.in0(_handshake_cond_br13_outFalse),
		.in0_valid(_handshake_cond_br13_outFalse_valid),
		.in0_ready(_handshake_sink7_in0_ready)
	);
	handshake_cond_br_in_ui1_2ins_2outs_ctrl handshake_cond_br14(
		.cond(_handshake_buffer97_out0),
		.cond_valid(_handshake_buffer97_out0_valid),
		.data_valid(_handshake_buffer79_out0_valid),
		.outTrue_ready(_handshake_buffer120_in0_ready),
		.outFalse_ready(_handshake_buffer119_in0_ready),
		.cond_ready(_handshake_cond_br14_cond_ready),
		.data_ready(_handshake_cond_br14_data_ready),
		.outTrue_valid(_handshake_cond_br14_outTrue_valid),
		.outFalse_valid(_handshake_cond_br14_outFalse_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer119(
		.in0_valid(_handshake_cond_br14_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux0_in1_ready),
		.in0_ready(_handshake_buffer119_in0_ready),
		.out0_valid(_handshake_buffer119_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer120(
		.in0_valid(_handshake_cond_br14_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork17_in0_ready),
		.in0_ready(_handshake_buffer120_in0_ready),
		.out0_valid(_handshake_buffer120_out0_valid)
	);
	handshake_fork_1ins_6outs_ctrl handshake_fork17(
		.in0_valid(_handshake_buffer120_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer126_in0_ready),
		.out1_ready(_handshake_buffer125_in0_ready),
		.out2_ready(_handshake_buffer124_in0_ready),
		.out3_ready(_handshake_buffer123_in0_ready),
		.out4_ready(_handshake_buffer122_in0_ready),
		.out5_ready(_handshake_buffer121_in0_ready),
		.in0_ready(_handshake_fork17_in0_ready),
		.out0_valid(_handshake_fork17_out0_valid),
		.out1_valid(_handshake_fork17_out1_valid),
		.out2_valid(_handshake_fork17_out2_valid),
		.out3_valid(_handshake_fork17_out3_valid),
		.out4_valid(_handshake_fork17_out4_valid),
		.out5_valid(_handshake_fork17_out5_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer121(
		.in0_valid(_handshake_fork17_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant6_ctrl_ready),
		.in0_ready(_handshake_buffer121_in0_ready),
		.out0_valid(_handshake_buffer121_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer122(
		.in0_valid(_handshake_fork17_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant7_ctrl_ready),
		.in0_ready(_handshake_buffer122_in0_ready),
		.out0_valid(_handshake_buffer122_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer123(
		.in0_valid(_handshake_fork17_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant8_ctrl_ready),
		.in0_ready(_handshake_buffer123_in0_ready),
		.out0_valid(_handshake_buffer123_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer124(
		.in0_valid(_handshake_fork17_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant9_ctrl_ready),
		.in0_ready(_handshake_buffer124_in0_ready),
		.out0_valid(_handshake_buffer124_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer125(
		.in0_valid(_handshake_fork17_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join3_in0_ready),
		.in0_ready(_handshake_buffer125_in0_ready),
		.out0_valid(_handshake_buffer125_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer126(
		.in0_valid(_handshake_fork17_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load0_ctrl_ready),
		.in0_ready(_handshake_buffer126_in0_ready),
		.out0_valid(_handshake_buffer126_out0_valid)
	);
	handshake_join_2ins_1outs_ctrl handshake_join3(
		.in0_valid(_handshake_buffer125_out0_valid),
		.in1_valid(_handshake_buffer13_out0_valid),
		.out0_ready(_handshake_buffer127_in0_ready),
		.in0_ready(_handshake_join3_in0_ready),
		.in1_ready(_handshake_join3_in1_ready),
		.out0_valid(_handshake_join3_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer127(
		.in0_valid(_handshake_join3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_control_merge1_in0_ready),
		.in0_ready(_handshake_buffer127_in0_ready),
		.out0_valid(_handshake_buffer127_out0_valid)
	);
	handshake_constant_c30_out_ui64 handshake_constant6(
		.ctrl_valid(_handshake_buffer121_out0_valid),
		.out0_ready(_handshake_buffer128_in0_ready),
		.ctrl_ready(_handshake_constant6_ctrl_ready),
		.out0(_handshake_constant6_out0),
		.out0_valid(_handshake_constant6_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer128(
		.in0(_handshake_constant6_out0),
		.in0_valid(_handshake_constant6_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli0_in1_ready),
		.in0_ready(_handshake_buffer128_in0_ready),
		.out0(_handshake_buffer128_out0),
		.out0_valid(_handshake_buffer128_out0_valid)
	);
	arith_muli_in_ui64_ui64_out_ui64 arith_muli0(
		.in0(_handshake_buffer115_out0),
		.in0_valid(_handshake_buffer115_out0_valid),
		.in1(_handshake_buffer128_out0),
		.in1_valid(_handshake_buffer128_out0_valid),
		.out0_ready(_handshake_buffer129_in0_ready),
		.in0_ready(_arith_muli0_in0_ready),
		.in1_ready(_arith_muli0_in1_ready),
		.out0(_arith_muli0_out0),
		.out0_valid(_arith_muli0_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer129(
		.in0(_arith_muli0_out0),
		.in0_valid(_arith_muli0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi0_in0_ready),
		.in0_ready(_handshake_buffer129_in0_ready),
		.out0(_handshake_buffer129_out0),
		.out0_valid(_handshake_buffer129_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi0(
		.in0(_handshake_buffer129_out0),
		.in0_valid(_handshake_buffer129_out0_valid),
		.in1(_handshake_buffer99_out0),
		.in1_valid(_handshake_buffer99_out0_valid),
		.out0_ready(_handshake_buffer130_in0_ready),
		.in0_ready(_arith_addi0_in0_ready),
		.in1_ready(_arith_addi0_in1_ready),
		.out0(_arith_addi0_out0),
		.out0_valid(_arith_addi0_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer130(
		.in0(_arith_addi0_out0),
		.in0_valid(_arith_addi0_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load0_addrIn0_ready),
		.in0_ready(_handshake_buffer130_in0_ready),
		.out0(_handshake_buffer130_out0),
		.out0_valid(_handshake_buffer130_out0_valid)
	);
	handshake_load_in_ui64_ui32_out_ui32_ui64 handshake_load0(
		.addrIn0(_handshake_buffer130_out0),
		.addrIn0_valid(_handshake_buffer130_out0_valid),
		.dataFromMem(_handshake_buffer12_out0),
		.dataFromMem_valid(_handshake_buffer12_out0_valid),
		.ctrl_valid(_handshake_buffer126_out0_valid),
		.dataOut_ready(_handshake_buffer132_in0_ready),
		.addrOut0_ready(_handshake_buffer131_in0_ready),
		.addrIn0_ready(_handshake_load0_addrIn0_ready),
		.dataFromMem_ready(_handshake_load0_dataFromMem_ready),
		.ctrl_ready(_handshake_load0_ctrl_ready),
		.dataOut(_handshake_load0_dataOut),
		.dataOut_valid(_handshake_load0_dataOut_valid),
		.addrOut0(_handshake_load0_addrOut0),
		.addrOut0_valid(_handshake_load0_addrOut0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer131(
		.in0(_handshake_load0_addrOut0),
		.in0_valid(_handshake_load0_addrOut0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_index_cast0_in0_ready),
		.in0_ready(_handshake_buffer131_in0_ready),
		.out0(_handshake_buffer131_out0),
		.out0_valid(_handshake_buffer131_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer132(
		.in0(_handshake_load0_dataOut),
		.in0_valid(_handshake_load0_dataOut_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli1_in0_ready),
		.in0_ready(_handshake_buffer132_in0_ready),
		.out0(_handshake_buffer132_out0),
		.out0_valid(_handshake_buffer132_out0_valid)
	);
	arith_muli_in_ui32_ui32_out_ui32 arith_muli1(
		.in0(_handshake_buffer132_out0),
		.in0_valid(_handshake_buffer132_out0_valid),
		.in1(_handshake_buffer105_out0),
		.in1_valid(_handshake_buffer105_out0_valid),
		.out0_ready(_handshake_buffer133_in0_ready),
		.in0_ready(_arith_muli1_in0_ready),
		.in1_ready(_arith_muli1_in1_ready),
		.out0(_arith_muli1_out0),
		.out0_valid(_arith_muli1_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer133(
		.in0(_arith_muli1_out0),
		.in0_valid(_arith_muli1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux15_in0_ready),
		.in0_ready(_handshake_buffer133_in0_ready),
		.out0(_handshake_buffer133_out0),
		.out0_valid(_handshake_buffer133_out0_valid)
	);
	handshake_constant_c0_out_ui64 handshake_constant7(
		.ctrl_valid(_handshake_buffer122_out0_valid),
		.out0_ready(_handshake_buffer134_in0_ready),
		.ctrl_ready(_handshake_constant7_ctrl_ready),
		.out0(_handshake_constant7_out0),
		.out0_valid(_handshake_constant7_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer134(
		.in0(_handshake_constant7_out0),
		.in0_valid(_handshake_constant7_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux14_in0_ready),
		.in0_ready(_handshake_buffer134_in0_ready),
		.out0(_handshake_buffer134_out0),
		.out0_valid(_handshake_buffer134_out0_valid)
	);
	handshake_constant_c20_out_ui64 handshake_constant8(
		.ctrl_valid(_handshake_buffer123_out0_valid),
		.out0_ready(_handshake_buffer135_in0_ready),
		.ctrl_ready(_handshake_constant8_ctrl_ready),
		.out0(_handshake_constant8_out0),
		.out0_valid(_handshake_constant8_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer135(
		.in0(_handshake_constant8_out0),
		.in0_valid(_handshake_constant8_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux24_in0_ready),
		.in0_ready(_handshake_buffer135_in0_ready),
		.out0(_handshake_buffer135_out0),
		.out0_valid(_handshake_buffer135_out0_valid)
	);
	handshake_constant_c1_out_ui64 handshake_constant9(
		.ctrl_valid(_handshake_buffer124_out0_valid),
		.out0_ready(_handshake_buffer136_in0_ready),
		.ctrl_ready(_handshake_constant9_ctrl_ready),
		.out0(_handshake_constant9_out0),
		.out0_valid(_handshake_constant9_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer136(
		.in0(_handshake_constant9_out0),
		.in0_valid(_handshake_constant9_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux25_in0_ready),
		.in0_ready(_handshake_buffer136_in0_ready),
		.out0(_handshake_buffer136_out0),
		.out0_valid(_handshake_buffer136_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux14(
		.select(_handshake_buffer155_out0),
		.select_valid(_handshake_buffer155_out0_valid),
		.in0(_handshake_buffer134_out0),
		.in0_valid(_handshake_buffer134_out0_valid),
		.in1(_handshake_buffer243_out0),
		.in1_valid(_handshake_buffer243_out0_valid),
		.out0_ready(_handshake_buffer137_in0_ready),
		.select_ready(_handshake_mux14_select_ready),
		.in0_ready(_handshake_mux14_in0_ready),
		.in1_ready(_handshake_mux14_in1_ready),
		.out0(_handshake_mux14_out0),
		.out0_valid(_handshake_mux14_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer137(
		.in0(_handshake_mux14_out0),
		.in0_valid(_handshake_mux14_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork18_in0_ready),
		.in0_ready(_handshake_buffer137_in0_ready),
		.out0(_handshake_buffer137_out0),
		.out0_valid(_handshake_buffer137_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork18(
		.in0(_handshake_buffer137_out0),
		.in0_valid(_handshake_buffer137_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer139_in0_ready),
		.out1_ready(_handshake_buffer138_in0_ready),
		.in0_ready(_handshake_fork18_in0_ready),
		.out0(_handshake_fork18_out0),
		.out0_valid(_handshake_fork18_out0_valid),
		.out1(_handshake_fork18_out1),
		.out1_valid(_handshake_fork18_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer138(
		.in0(_handshake_fork18_out1),
		.in0_valid(_handshake_fork18_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi2_in0_ready),
		.in0_ready(_handshake_buffer138_in0_ready),
		.out0(_handshake_buffer138_out0),
		.out0_valid(_handshake_buffer138_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer139(
		.in0(_handshake_fork18_out0),
		.in0_valid(_handshake_fork18_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br15_data_ready),
		.in0_ready(_handshake_buffer139_in0_ready),
		.out0(_handshake_buffer139_out0),
		.out0_valid(_handshake_buffer139_out0_valid)
	);
	handshake_mux_in_ui64_ui32_ui32_out_ui32 handshake_mux15(
		.select(_handshake_buffer156_out0),
		.select_valid(_handshake_buffer156_out0_valid),
		.in0(_handshake_buffer133_out0),
		.in0_valid(_handshake_buffer133_out0_valid),
		.in1(_handshake_buffer242_out0),
		.in1_valid(_handshake_buffer242_out0_valid),
		.out0_ready(_handshake_buffer140_in0_ready),
		.select_ready(_handshake_mux15_select_ready),
		.in0_ready(_handshake_mux15_in0_ready),
		.in1_ready(_handshake_mux15_in1_ready),
		.out0(_handshake_mux15_out0),
		.out0_valid(_handshake_mux15_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer140(
		.in0(_handshake_mux15_out0),
		.in0_valid(_handshake_mux15_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br16_data_ready),
		.in0_ready(_handshake_buffer140_in0_ready),
		.out0(_handshake_buffer140_out0),
		.out0_valid(_handshake_buffer140_out0_valid)
	);
	handshake_mux_in_ui64_ui32_ui32_out_ui32 handshake_mux16(
		.select(_handshake_buffer157_out0),
		.select_valid(_handshake_buffer157_out0_valid),
		.in0(_handshake_buffer102_out0),
		.in0_valid(_handshake_buffer102_out0_valid),
		.in1(_handshake_buffer190_out0),
		.in1_valid(_handshake_buffer190_out0_valid),
		.out0_ready(_handshake_buffer141_in0_ready),
		.select_ready(_handshake_mux16_select_ready),
		.in0_ready(_handshake_mux16_in0_ready),
		.in1_ready(_handshake_mux16_in1_ready),
		.out0(_handshake_mux16_out0),
		.out0_valid(_handshake_mux16_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer141(
		.in0(_handshake_mux16_out0),
		.in0_valid(_handshake_mux16_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br17_data_ready),
		.in0_ready(_handshake_buffer141_in0_ready),
		.out0(_handshake_buffer141_out0),
		.out0_valid(_handshake_buffer141_out0_valid)
	);
	handshake_mux_in_ui64_ui32_ui32_out_ui32 handshake_mux17(
		.select(_handshake_buffer158_out0),
		.select_valid(_handshake_buffer158_out0_valid),
		.in0(_handshake_buffer106_out0),
		.in0_valid(_handshake_buffer106_out0_valid),
		.in1(_handshake_buffer192_out0),
		.in1_valid(_handshake_buffer192_out0_valid),
		.out0_ready(_handshake_buffer142_in0_ready),
		.select_ready(_handshake_mux17_select_ready),
		.in0_ready(_handshake_mux17_in0_ready),
		.in1_ready(_handshake_mux17_in1_ready),
		.out0(_handshake_mux17_out0),
		.out0_valid(_handshake_mux17_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer142(
		.in0(_handshake_mux17_out0),
		.in0_valid(_handshake_mux17_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br18_data_ready),
		.in0_ready(_handshake_buffer142_in0_ready),
		.out0(_handshake_buffer142_out0),
		.out0_valid(_handshake_buffer142_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux18(
		.select(_handshake_buffer159_out0),
		.select_valid(_handshake_buffer159_out0_valid),
		.in0(_handshake_buffer108_out0),
		.in0_valid(_handshake_buffer108_out0_valid),
		.in1(_handshake_buffer194_out0),
		.in1_valid(_handshake_buffer194_out0_valid),
		.out0_ready(_handshake_buffer143_in0_ready),
		.select_ready(_handshake_mux18_select_ready),
		.in0_ready(_handshake_mux18_in0_ready),
		.in1_ready(_handshake_mux18_in1_ready),
		.out0(_handshake_mux18_out0),
		.out0_valid(_handshake_mux18_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer143(
		.in0(_handshake_mux18_out0),
		.in0_valid(_handshake_mux18_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br19_data_ready),
		.in0_ready(_handshake_buffer143_in0_ready),
		.out0(_handshake_buffer143_out0),
		.out0_valid(_handshake_buffer143_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux19(
		.select(_handshake_buffer160_out0),
		.select_valid(_handshake_buffer160_out0_valid),
		.in0(_handshake_buffer110_out0),
		.in0_valid(_handshake_buffer110_out0_valid),
		.in1(_handshake_buffer196_out0),
		.in1_valid(_handshake_buffer196_out0_valid),
		.out0_ready(_handshake_buffer144_in0_ready),
		.select_ready(_handshake_mux19_select_ready),
		.in0_ready(_handshake_mux19_in0_ready),
		.in1_ready(_handshake_mux19_in1_ready),
		.out0(_handshake_mux19_out0),
		.out0_valid(_handshake_mux19_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer144(
		.in0(_handshake_mux19_out0),
		.in0_valid(_handshake_mux19_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br20_data_ready),
		.in0_ready(_handshake_buffer144_in0_ready),
		.out0(_handshake_buffer144_out0),
		.out0_valid(_handshake_buffer144_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux20(
		.select(_handshake_buffer161_out0),
		.select_valid(_handshake_buffer161_out0_valid),
		.in0(_handshake_buffer116_out0),
		.in0_valid(_handshake_buffer116_out0_valid),
		.in1(_handshake_buffer202_out0),
		.in1_valid(_handshake_buffer202_out0_valid),
		.out0_ready(_handshake_buffer145_in0_ready),
		.select_ready(_handshake_mux20_select_ready),
		.in0_ready(_handshake_mux20_in0_ready),
		.in1_ready(_handshake_mux20_in1_ready),
		.out0(_handshake_mux20_out0),
		.out0_valid(_handshake_mux20_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer145(
		.in0(_handshake_mux20_out0),
		.in0_valid(_handshake_mux20_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br21_data_ready),
		.in0_ready(_handshake_buffer145_in0_ready),
		.out0(_handshake_buffer145_out0),
		.out0_valid(_handshake_buffer145_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux21(
		.select(_handshake_buffer162_out0),
		.select_valid(_handshake_buffer162_out0_valid),
		.in0(_handshake_buffer117_out0),
		.in0_valid(_handshake_buffer117_out0_valid),
		.in1(_handshake_buffer204_out0),
		.in1_valid(_handshake_buffer204_out0_valid),
		.out0_ready(_handshake_buffer146_in0_ready),
		.select_ready(_handshake_mux21_select_ready),
		.in0_ready(_handshake_mux21_in0_ready),
		.in1_ready(_handshake_mux21_in1_ready),
		.out0(_handshake_mux21_out0),
		.out0_valid(_handshake_mux21_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer146(
		.in0(_handshake_mux21_out0),
		.in0_valid(_handshake_mux21_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br22_data_ready),
		.in0_ready(_handshake_buffer146_in0_ready),
		.out0(_handshake_buffer146_out0),
		.out0_valid(_handshake_buffer146_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux22(
		.select(_handshake_buffer163_out0),
		.select_valid(_handshake_buffer163_out0_valid),
		.in0(_handshake_buffer118_out0),
		.in0_valid(_handshake_buffer118_out0_valid),
		.in1(_handshake_buffer206_out0),
		.in1_valid(_handshake_buffer206_out0_valid),
		.out0_ready(_handshake_buffer147_in0_ready),
		.select_ready(_handshake_mux22_select_ready),
		.in0_ready(_handshake_mux22_in0_ready),
		.in1_ready(_handshake_mux22_in1_ready),
		.out0(_handshake_mux22_out0),
		.out0_valid(_handshake_mux22_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer147(
		.in0(_handshake_mux22_out0),
		.in0_valid(_handshake_mux22_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br23_data_ready),
		.in0_ready(_handshake_buffer147_in0_ready),
		.out0(_handshake_buffer147_out0),
		.out0_valid(_handshake_buffer147_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux23(
		.select(_handshake_buffer164_out0),
		.select_valid(_handshake_buffer164_out0_valid),
		.in0(_handshake_buffer100_out0),
		.in0_valid(_handshake_buffer100_out0_valid),
		.in1(_handshake_buffer214_out0),
		.in1_valid(_handshake_buffer214_out0_valid),
		.out0_ready(_handshake_buffer148_in0_ready),
		.select_ready(_handshake_mux23_select_ready),
		.in0_ready(_handshake_mux23_in0_ready),
		.in1_ready(_handshake_mux23_in1_ready),
		.out0(_handshake_mux23_out0),
		.out0_valid(_handshake_mux23_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer148(
		.in0(_handshake_mux23_out0),
		.in0_valid(_handshake_mux23_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br24_data_ready),
		.in0_ready(_handshake_buffer148_in0_ready),
		.out0(_handshake_buffer148_out0),
		.out0_valid(_handshake_buffer148_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux24(
		.select(_handshake_buffer165_out0),
		.select_valid(_handshake_buffer165_out0_valid),
		.in0(_handshake_buffer135_out0),
		.in0_valid(_handshake_buffer135_out0_valid),
		.in1(_handshake_buffer215_out0),
		.in1_valid(_handshake_buffer215_out0_valid),
		.out0_ready(_handshake_buffer149_in0_ready),
		.select_ready(_handshake_mux24_select_ready),
		.in0_ready(_handshake_mux24_in0_ready),
		.in1_ready(_handshake_mux24_in1_ready),
		.out0(_handshake_mux24_out0),
		.out0_valid(_handshake_mux24_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer149(
		.in0(_handshake_mux24_out0),
		.in0_valid(_handshake_mux24_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork19_in0_ready),
		.in0_ready(_handshake_buffer149_in0_ready),
		.out0(_handshake_buffer149_out0),
		.out0_valid(_handshake_buffer149_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork19(
		.in0(_handshake_buffer149_out0),
		.in0_valid(_handshake_buffer149_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer151_in0_ready),
		.out1_ready(_handshake_buffer150_in0_ready),
		.in0_ready(_handshake_fork19_in0_ready),
		.out0(_handshake_fork19_out0),
		.out0_valid(_handshake_fork19_out0_valid),
		.out1(_handshake_fork19_out1),
		.out1_valid(_handshake_fork19_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer150(
		.in0(_handshake_fork19_out1),
		.in0_valid(_handshake_fork19_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_cmpi2_in1_ready),
		.in0_ready(_handshake_buffer150_in0_ready),
		.out0(_handshake_buffer150_out0),
		.out0_valid(_handshake_buffer150_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer151(
		.in0(_handshake_fork19_out0),
		.in0_valid(_handshake_fork19_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br25_data_ready),
		.in0_ready(_handshake_buffer151_in0_ready),
		.out0(_handshake_buffer151_out0),
		.out0_valid(_handshake_buffer151_out0_valid)
	);
	handshake_mux_in_ui64_ui64_ui64_out_ui64 handshake_mux25(
		.select(_handshake_buffer166_out0),
		.select_valid(_handshake_buffer166_out0_valid),
		.in0(_handshake_buffer136_out0),
		.in0_valid(_handshake_buffer136_out0_valid),
		.in1(_handshake_buffer218_out0),
		.in1_valid(_handshake_buffer218_out0_valid),
		.out0_ready(_handshake_buffer152_in0_ready),
		.select_ready(_handshake_mux25_select_ready),
		.in0_ready(_handshake_mux25_in0_ready),
		.in1_ready(_handshake_mux25_in1_ready),
		.out0(_handshake_mux25_out0),
		.out0_valid(_handshake_mux25_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer152(
		.in0(_handshake_mux25_out0),
		.in0_valid(_handshake_mux25_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br26_data_ready),
		.in0_ready(_handshake_buffer152_in0_ready),
		.out0(_handshake_buffer152_out0),
		.out0_valid(_handshake_buffer152_out0_valid)
	);
	handshake_control_merge_out_ui64_2ins_2outs_ctrl handshake_control_merge1(
		.in0_valid(_handshake_buffer127_out0_valid),
		.in1_valid(_handshake_buffer229_out0_valid),
		.clock(clock),
		.reset(reset),
		.dataOut_ready(_handshake_buffer154_in0_ready),
		.index_ready(_handshake_buffer153_in0_ready),
		.in0_ready(_handshake_control_merge1_in0_ready),
		.in1_ready(_handshake_control_merge1_in1_ready),
		.dataOut_valid(_handshake_control_merge1_dataOut_valid),
		.index(_handshake_control_merge1_index),
		.index_valid(_handshake_control_merge1_index_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer153(
		.in0(_handshake_control_merge1_index),
		.in0_valid(_handshake_control_merge1_index_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork20_in0_ready),
		.in0_ready(_handshake_buffer153_in0_ready),
		.out0(_handshake_buffer153_out0),
		.out0_valid(_handshake_buffer153_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer154(
		.in0_valid(_handshake_control_merge1_dataOut_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br27_data_ready),
		.in0_ready(_handshake_buffer154_in0_ready),
		.out0_valid(_handshake_buffer154_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64_ui64 handshake_fork20(
		.in0(_handshake_buffer153_out0),
		.in0_valid(_handshake_buffer153_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer166_in0_ready),
		.out1_ready(_handshake_buffer165_in0_ready),
		.out2_ready(_handshake_buffer164_in0_ready),
		.out3_ready(_handshake_buffer163_in0_ready),
		.out4_ready(_handshake_buffer162_in0_ready),
		.out5_ready(_handshake_buffer161_in0_ready),
		.out6_ready(_handshake_buffer160_in0_ready),
		.out7_ready(_handshake_buffer159_in0_ready),
		.out8_ready(_handshake_buffer158_in0_ready),
		.out9_ready(_handshake_buffer157_in0_ready),
		.out10_ready(_handshake_buffer156_in0_ready),
		.out11_ready(_handshake_buffer155_in0_ready),
		.in0_ready(_handshake_fork20_in0_ready),
		.out0(_handshake_fork20_out0),
		.out0_valid(_handshake_fork20_out0_valid),
		.out1(_handshake_fork20_out1),
		.out1_valid(_handshake_fork20_out1_valid),
		.out2(_handshake_fork20_out2),
		.out2_valid(_handshake_fork20_out2_valid),
		.out3(_handshake_fork20_out3),
		.out3_valid(_handshake_fork20_out3_valid),
		.out4(_handshake_fork20_out4),
		.out4_valid(_handshake_fork20_out4_valid),
		.out5(_handshake_fork20_out5),
		.out5_valid(_handshake_fork20_out5_valid),
		.out6(_handshake_fork20_out6),
		.out6_valid(_handshake_fork20_out6_valid),
		.out7(_handshake_fork20_out7),
		.out7_valid(_handshake_fork20_out7_valid),
		.out8(_handshake_fork20_out8),
		.out8_valid(_handshake_fork20_out8_valid),
		.out9(_handshake_fork20_out9),
		.out9_valid(_handshake_fork20_out9_valid),
		.out10(_handshake_fork20_out10),
		.out10_valid(_handshake_fork20_out10_valid),
		.out11(_handshake_fork20_out11),
		.out11_valid(_handshake_fork20_out11_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer155(
		.in0(_handshake_fork20_out11),
		.in0_valid(_handshake_fork20_out11_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux14_select_ready),
		.in0_ready(_handshake_buffer155_in0_ready),
		.out0(_handshake_buffer155_out0),
		.out0_valid(_handshake_buffer155_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer156(
		.in0(_handshake_fork20_out10),
		.in0_valid(_handshake_fork20_out10_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux15_select_ready),
		.in0_ready(_handshake_buffer156_in0_ready),
		.out0(_handshake_buffer156_out0),
		.out0_valid(_handshake_buffer156_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer157(
		.in0(_handshake_fork20_out9),
		.in0_valid(_handshake_fork20_out9_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux16_select_ready),
		.in0_ready(_handshake_buffer157_in0_ready),
		.out0(_handshake_buffer157_out0),
		.out0_valid(_handshake_buffer157_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer158(
		.in0(_handshake_fork20_out8),
		.in0_valid(_handshake_fork20_out8_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux17_select_ready),
		.in0_ready(_handshake_buffer158_in0_ready),
		.out0(_handshake_buffer158_out0),
		.out0_valid(_handshake_buffer158_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer159(
		.in0(_handshake_fork20_out7),
		.in0_valid(_handshake_fork20_out7_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux18_select_ready),
		.in0_ready(_handshake_buffer159_in0_ready),
		.out0(_handshake_buffer159_out0),
		.out0_valid(_handshake_buffer159_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer160(
		.in0(_handshake_fork20_out6),
		.in0_valid(_handshake_fork20_out6_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux19_select_ready),
		.in0_ready(_handshake_buffer160_in0_ready),
		.out0(_handshake_buffer160_out0),
		.out0_valid(_handshake_buffer160_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer161(
		.in0(_handshake_fork20_out5),
		.in0_valid(_handshake_fork20_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux20_select_ready),
		.in0_ready(_handshake_buffer161_in0_ready),
		.out0(_handshake_buffer161_out0),
		.out0_valid(_handshake_buffer161_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer162(
		.in0(_handshake_fork20_out4),
		.in0_valid(_handshake_fork20_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux21_select_ready),
		.in0_ready(_handshake_buffer162_in0_ready),
		.out0(_handshake_buffer162_out0),
		.out0_valid(_handshake_buffer162_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer163(
		.in0(_handshake_fork20_out3),
		.in0_valid(_handshake_fork20_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux22_select_ready),
		.in0_ready(_handshake_buffer163_in0_ready),
		.out0(_handshake_buffer163_out0),
		.out0_valid(_handshake_buffer163_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer164(
		.in0(_handshake_fork20_out2),
		.in0_valid(_handshake_fork20_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux23_select_ready),
		.in0_ready(_handshake_buffer164_in0_ready),
		.out0(_handshake_buffer164_out0),
		.out0_valid(_handshake_buffer164_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer165(
		.in0(_handshake_fork20_out1),
		.in0_valid(_handshake_fork20_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux24_select_ready),
		.in0_ready(_handshake_buffer165_in0_ready),
		.out0(_handshake_buffer165_out0),
		.out0_valid(_handshake_buffer165_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer166(
		.in0(_handshake_fork20_out0),
		.in0_valid(_handshake_fork20_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux25_select_ready),
		.in0_ready(_handshake_buffer166_in0_ready),
		.out0(_handshake_buffer166_out0),
		.out0_valid(_handshake_buffer166_out0_valid)
	);
	arith_cmpi_in_ui64_ui64_out_ui1_slt arith_cmpi2(
		.in0(_handshake_buffer138_out0),
		.in0_valid(_handshake_buffer138_out0_valid),
		.in1(_handshake_buffer150_out0),
		.in1_valid(_handshake_buffer150_out0_valid),
		.out0_ready(_handshake_buffer167_in0_ready),
		.in0_ready(_arith_cmpi2_in0_ready),
		.in1_ready(_arith_cmpi2_in1_ready),
		.out0(_arith_cmpi2_out0),
		.out0_valid(_arith_cmpi2_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer167(
		.in0(_arith_cmpi2_out0),
		.in0_valid(_arith_cmpi2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork21_in0_ready),
		.in0_ready(_handshake_buffer167_in0_ready),
		.out0(_handshake_buffer167_out0),
		.out0_valid(_handshake_buffer167_out0_valid)
	);
	handshake_fork_in_ui1_out_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1_ui1 handshake_fork21(
		.in0(_handshake_buffer167_out0),
		.in0_valid(_handshake_buffer167_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer180_in0_ready),
		.out1_ready(_handshake_buffer179_in0_ready),
		.out2_ready(_handshake_buffer178_in0_ready),
		.out3_ready(_handshake_buffer177_in0_ready),
		.out4_ready(_handshake_buffer176_in0_ready),
		.out5_ready(_handshake_buffer175_in0_ready),
		.out6_ready(_handshake_buffer174_in0_ready),
		.out7_ready(_handshake_buffer173_in0_ready),
		.out8_ready(_handshake_buffer172_in0_ready),
		.out9_ready(_handshake_buffer171_in0_ready),
		.out10_ready(_handshake_buffer170_in0_ready),
		.out11_ready(_handshake_buffer169_in0_ready),
		.out12_ready(_handshake_buffer168_in0_ready),
		.in0_ready(_handshake_fork21_in0_ready),
		.out0(_handshake_fork21_out0),
		.out0_valid(_handshake_fork21_out0_valid),
		.out1(_handshake_fork21_out1),
		.out1_valid(_handshake_fork21_out1_valid),
		.out2(_handshake_fork21_out2),
		.out2_valid(_handshake_fork21_out2_valid),
		.out3(_handshake_fork21_out3),
		.out3_valid(_handshake_fork21_out3_valid),
		.out4(_handshake_fork21_out4),
		.out4_valid(_handshake_fork21_out4_valid),
		.out5(_handshake_fork21_out5),
		.out5_valid(_handshake_fork21_out5_valid),
		.out6(_handshake_fork21_out6),
		.out6_valid(_handshake_fork21_out6_valid),
		.out7(_handshake_fork21_out7),
		.out7_valid(_handshake_fork21_out7_valid),
		.out8(_handshake_fork21_out8),
		.out8_valid(_handshake_fork21_out8_valid),
		.out9(_handshake_fork21_out9),
		.out9_valid(_handshake_fork21_out9_valid),
		.out10(_handshake_fork21_out10),
		.out10_valid(_handshake_fork21_out10_valid),
		.out11(_handshake_fork21_out11),
		.out11_valid(_handshake_fork21_out11_valid),
		.out12(_handshake_fork21_out12),
		.out12_valid(_handshake_fork21_out12_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer168(
		.in0(_handshake_fork21_out12),
		.in0_valid(_handshake_fork21_out12_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br15_cond_ready),
		.in0_ready(_handshake_buffer168_in0_ready),
		.out0(_handshake_buffer168_out0),
		.out0_valid(_handshake_buffer168_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer169(
		.in0(_handshake_fork21_out11),
		.in0_valid(_handshake_fork21_out11_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br16_cond_ready),
		.in0_ready(_handshake_buffer169_in0_ready),
		.out0(_handshake_buffer169_out0),
		.out0_valid(_handshake_buffer169_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer170(
		.in0(_handshake_fork21_out10),
		.in0_valid(_handshake_fork21_out10_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br17_cond_ready),
		.in0_ready(_handshake_buffer170_in0_ready),
		.out0(_handshake_buffer170_out0),
		.out0_valid(_handshake_buffer170_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer171(
		.in0(_handshake_fork21_out9),
		.in0_valid(_handshake_fork21_out9_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br18_cond_ready),
		.in0_ready(_handshake_buffer171_in0_ready),
		.out0(_handshake_buffer171_out0),
		.out0_valid(_handshake_buffer171_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer172(
		.in0(_handshake_fork21_out8),
		.in0_valid(_handshake_fork21_out8_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br19_cond_ready),
		.in0_ready(_handshake_buffer172_in0_ready),
		.out0(_handshake_buffer172_out0),
		.out0_valid(_handshake_buffer172_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer173(
		.in0(_handshake_fork21_out7),
		.in0_valid(_handshake_fork21_out7_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br20_cond_ready),
		.in0_ready(_handshake_buffer173_in0_ready),
		.out0(_handshake_buffer173_out0),
		.out0_valid(_handshake_buffer173_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer174(
		.in0(_handshake_fork21_out6),
		.in0_valid(_handshake_fork21_out6_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br21_cond_ready),
		.in0_ready(_handshake_buffer174_in0_ready),
		.out0(_handshake_buffer174_out0),
		.out0_valid(_handshake_buffer174_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer175(
		.in0(_handshake_fork21_out5),
		.in0_valid(_handshake_fork21_out5_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br22_cond_ready),
		.in0_ready(_handshake_buffer175_in0_ready),
		.out0(_handshake_buffer175_out0),
		.out0_valid(_handshake_buffer175_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer176(
		.in0(_handshake_fork21_out4),
		.in0_valid(_handshake_fork21_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br23_cond_ready),
		.in0_ready(_handshake_buffer176_in0_ready),
		.out0(_handshake_buffer176_out0),
		.out0_valid(_handshake_buffer176_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer177(
		.in0(_handshake_fork21_out3),
		.in0_valid(_handshake_fork21_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br24_cond_ready),
		.in0_ready(_handshake_buffer177_in0_ready),
		.out0(_handshake_buffer177_out0),
		.out0_valid(_handshake_buffer177_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer178(
		.in0(_handshake_fork21_out2),
		.in0_valid(_handshake_fork21_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br25_cond_ready),
		.in0_ready(_handshake_buffer178_in0_ready),
		.out0(_handshake_buffer178_out0),
		.out0_valid(_handshake_buffer178_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer179(
		.in0(_handshake_fork21_out1),
		.in0_valid(_handshake_fork21_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br26_cond_ready),
		.in0_ready(_handshake_buffer179_in0_ready),
		.out0(_handshake_buffer179_out0),
		.out0_valid(_handshake_buffer179_out0_valid)
	);
	handshake_buffer_in_ui1_out_ui1_2slots_seq handshake_buffer180(
		.in0(_handshake_fork21_out0),
		.in0_valid(_handshake_fork21_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_cond_br27_cond_ready),
		.in0_ready(_handshake_buffer180_in0_ready),
		.out0(_handshake_buffer180_out0),
		.out0_valid(_handshake_buffer180_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br15(
		.cond(_handshake_buffer168_out0),
		.cond_valid(_handshake_buffer168_out0_valid),
		.data(_handshake_buffer139_out0),
		.data_valid(_handshake_buffer139_out0_valid),
		.outTrue_ready(_handshake_buffer181_in0_ready),
		.outFalse_ready(_handshake_sink8_in0_ready),
		.cond_ready(_handshake_cond_br15_cond_ready),
		.data_ready(_handshake_cond_br15_data_ready),
		.outTrue(_handshake_cond_br15_outTrue),
		.outTrue_valid(_handshake_cond_br15_outTrue_valid),
		.outFalse(_handshake_cond_br15_outFalse),
		.outFalse_valid(_handshake_cond_br15_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer181(
		.in0(_handshake_cond_br15_outTrue),
		.in0_valid(_handshake_cond_br15_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork22_in0_ready),
		.in0_ready(_handshake_buffer181_in0_ready),
		.out0(_handshake_buffer181_out0),
		.out0_valid(_handshake_buffer181_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink8(
		.in0(_handshake_cond_br15_outFalse),
		.in0_valid(_handshake_cond_br15_outFalse_valid),
		.in0_ready(_handshake_sink8_in0_ready)
	);
	handshake_fork_in_ui64_out_ui64_ui64_ui64 handshake_fork22(
		.in0(_handshake_buffer181_out0),
		.in0_valid(_handshake_buffer181_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer184_in0_ready),
		.out1_ready(_handshake_buffer183_in0_ready),
		.out2_ready(_handshake_buffer182_in0_ready),
		.in0_ready(_handshake_fork22_in0_ready),
		.out0(_handshake_fork22_out0),
		.out0_valid(_handshake_fork22_out0_valid),
		.out1(_handshake_fork22_out1),
		.out1_valid(_handshake_fork22_out1_valid),
		.out2(_handshake_fork22_out2),
		.out2_valid(_handshake_fork22_out2_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer182(
		.in0(_handshake_fork22_out2),
		.in0_valid(_handshake_fork22_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi4_in0_ready),
		.in0_ready(_handshake_buffer182_in0_ready),
		.out0(_handshake_buffer182_out0),
		.out0_valid(_handshake_buffer182_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer183(
		.in0(_handshake_fork22_out1),
		.in0_valid(_handshake_fork22_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli4_in0_ready),
		.in0_ready(_handshake_buffer183_in0_ready),
		.out0(_handshake_buffer183_out0),
		.out0_valid(_handshake_buffer183_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer184(
		.in0(_handshake_fork22_out0),
		.in0_valid(_handshake_fork22_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi1_in1_ready),
		.in0_ready(_handshake_buffer184_in0_ready),
		.out0(_handshake_buffer184_out0),
		.out0_valid(_handshake_buffer184_out0_valid)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br16(
		.cond(_handshake_buffer169_out0),
		.cond_valid(_handshake_buffer169_out0_valid),
		.data(_handshake_buffer140_out0),
		.data_valid(_handshake_buffer140_out0_valid),
		.outTrue_ready(_handshake_buffer186_in0_ready),
		.outFalse_ready(_handshake_buffer185_in0_ready),
		.cond_ready(_handshake_cond_br16_cond_ready),
		.data_ready(_handshake_cond_br16_data_ready),
		.outTrue(_handshake_cond_br16_outTrue),
		.outTrue_valid(_handshake_cond_br16_outTrue_valid),
		.outFalse(_handshake_cond_br16_outFalse),
		.outFalse_valid(_handshake_cond_br16_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer185(
		.in0(_handshake_cond_br16_outFalse),
		.in0_valid(_handshake_cond_br16_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_store0_dataIn_ready),
		.in0_ready(_handshake_buffer185_in0_ready),
		.out0(_handshake_buffer185_out0),
		.out0_valid(_handshake_buffer185_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer186(
		.in0(_handshake_cond_br16_outTrue),
		.in0_valid(_handshake_cond_br16_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi3_in0_ready),
		.in0_ready(_handshake_buffer186_in0_ready),
		.out0(_handshake_buffer186_out0),
		.out0_valid(_handshake_buffer186_out0_valid)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br17(
		.cond(_handshake_buffer170_out0),
		.cond_valid(_handshake_buffer170_out0_valid),
		.data(_handshake_buffer141_out0),
		.data_valid(_handshake_buffer141_out0_valid),
		.outTrue_ready(_handshake_buffer188_in0_ready),
		.outFalse_ready(_handshake_buffer187_in0_ready),
		.cond_ready(_handshake_cond_br17_cond_ready),
		.data_ready(_handshake_cond_br17_data_ready),
		.outTrue(_handshake_cond_br17_outTrue),
		.outTrue_valid(_handshake_cond_br17_outTrue_valid),
		.outFalse(_handshake_cond_br17_outFalse),
		.outFalse_valid(_handshake_cond_br17_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer187(
		.in0(_handshake_cond_br17_outFalse),
		.in0_valid(_handshake_cond_br17_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux7_in1_ready),
		.in0_ready(_handshake_buffer187_in0_ready),
		.out0(_handshake_buffer187_out0),
		.out0_valid(_handshake_buffer187_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer188(
		.in0(_handshake_cond_br17_outTrue),
		.in0_valid(_handshake_cond_br17_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork23_in0_ready),
		.in0_ready(_handshake_buffer188_in0_ready),
		.out0(_handshake_buffer188_out0),
		.out0_valid(_handshake_buffer188_out0_valid)
	);
	handshake_fork_in_ui32_out_ui32_ui32 handshake_fork23(
		.in0(_handshake_buffer188_out0),
		.in0_valid(_handshake_buffer188_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer190_in0_ready),
		.out1_ready(_handshake_buffer189_in0_ready),
		.in0_ready(_handshake_fork23_in0_ready),
		.out0(_handshake_fork23_out0),
		.out0_valid(_handshake_fork23_out0_valid),
		.out1(_handshake_fork23_out1),
		.out1_valid(_handshake_fork23_out1_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer189(
		.in0(_handshake_fork23_out1),
		.in0_valid(_handshake_fork23_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli3_in0_ready),
		.in0_ready(_handshake_buffer189_in0_ready),
		.out0(_handshake_buffer189_out0),
		.out0_valid(_handshake_buffer189_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer190(
		.in0(_handshake_fork23_out0),
		.in0_valid(_handshake_fork23_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux16_in1_ready),
		.in0_ready(_handshake_buffer190_in0_ready),
		.out0(_handshake_buffer190_out0),
		.out0_valid(_handshake_buffer190_out0_valid)
	);
	handshake_cond_br_in_ui1_ui32_out_ui32_ui32 handshake_cond_br18(
		.cond(_handshake_buffer171_out0),
		.cond_valid(_handshake_buffer171_out0_valid),
		.data(_handshake_buffer142_out0),
		.data_valid(_handshake_buffer142_out0_valid),
		.outTrue_ready(_handshake_buffer192_in0_ready),
		.outFalse_ready(_handshake_buffer191_in0_ready),
		.cond_ready(_handshake_cond_br18_cond_ready),
		.data_ready(_handshake_cond_br18_data_ready),
		.outTrue(_handshake_cond_br18_outTrue),
		.outTrue_valid(_handshake_cond_br18_outTrue_valid),
		.outFalse(_handshake_cond_br18_outFalse),
		.outFalse_valid(_handshake_cond_br18_outFalse_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer191(
		.in0(_handshake_cond_br18_outFalse),
		.in0_valid(_handshake_cond_br18_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux8_in1_ready),
		.in0_ready(_handshake_buffer191_in0_ready),
		.out0(_handshake_buffer191_out0),
		.out0_valid(_handshake_buffer191_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer192(
		.in0(_handshake_cond_br18_outTrue),
		.in0_valid(_handshake_cond_br18_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux17_in1_ready),
		.in0_ready(_handshake_buffer192_in0_ready),
		.out0(_handshake_buffer192_out0),
		.out0_valid(_handshake_buffer192_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br19(
		.cond(_handshake_buffer172_out0),
		.cond_valid(_handshake_buffer172_out0_valid),
		.data(_handshake_buffer143_out0),
		.data_valid(_handshake_buffer143_out0_valid),
		.outTrue_ready(_handshake_buffer194_in0_ready),
		.outFalse_ready(_handshake_buffer193_in0_ready),
		.cond_ready(_handshake_cond_br19_cond_ready),
		.data_ready(_handshake_cond_br19_data_ready),
		.outTrue(_handshake_cond_br19_outTrue),
		.outTrue_valid(_handshake_cond_br19_outTrue_valid),
		.outFalse(_handshake_cond_br19_outFalse),
		.outFalse_valid(_handshake_cond_br19_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer193(
		.in0(_handshake_cond_br19_outFalse),
		.in0_valid(_handshake_cond_br19_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux9_in1_ready),
		.in0_ready(_handshake_buffer193_in0_ready),
		.out0(_handshake_buffer193_out0),
		.out0_valid(_handshake_buffer193_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer194(
		.in0(_handshake_cond_br19_outTrue),
		.in0_valid(_handshake_cond_br19_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux18_in1_ready),
		.in0_ready(_handshake_buffer194_in0_ready),
		.out0(_handshake_buffer194_out0),
		.out0_valid(_handshake_buffer194_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br20(
		.cond(_handshake_buffer173_out0),
		.cond_valid(_handshake_buffer173_out0_valid),
		.data(_handshake_buffer144_out0),
		.data_valid(_handshake_buffer144_out0_valid),
		.outTrue_ready(_handshake_buffer196_in0_ready),
		.outFalse_ready(_handshake_buffer195_in0_ready),
		.cond_ready(_handshake_cond_br20_cond_ready),
		.data_ready(_handshake_cond_br20_data_ready),
		.outTrue(_handshake_cond_br20_outTrue),
		.outTrue_valid(_handshake_cond_br20_outTrue_valid),
		.outFalse(_handshake_cond_br20_outFalse),
		.outFalse_valid(_handshake_cond_br20_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer195(
		.in0(_handshake_cond_br20_outFalse),
		.in0_valid(_handshake_cond_br20_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux10_in1_ready),
		.in0_ready(_handshake_buffer195_in0_ready),
		.out0(_handshake_buffer195_out0),
		.out0_valid(_handshake_buffer195_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer196(
		.in0(_handshake_cond_br20_outTrue),
		.in0_valid(_handshake_cond_br20_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux19_in1_ready),
		.in0_ready(_handshake_buffer196_in0_ready),
		.out0(_handshake_buffer196_out0),
		.out0_valid(_handshake_buffer196_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br21(
		.cond(_handshake_buffer174_out0),
		.cond_valid(_handshake_buffer174_out0_valid),
		.data(_handshake_buffer145_out0),
		.data_valid(_handshake_buffer145_out0_valid),
		.outTrue_ready(_handshake_buffer198_in0_ready),
		.outFalse_ready(_handshake_buffer197_in0_ready),
		.cond_ready(_handshake_cond_br21_cond_ready),
		.data_ready(_handshake_cond_br21_data_ready),
		.outTrue(_handshake_cond_br21_outTrue),
		.outTrue_valid(_handshake_cond_br21_outTrue_valid),
		.outFalse(_handshake_cond_br21_outFalse),
		.outFalse_valid(_handshake_cond_br21_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer197(
		.in0(_handshake_cond_br21_outFalse),
		.in0_valid(_handshake_cond_br21_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork24_in0_ready),
		.in0_ready(_handshake_buffer197_in0_ready),
		.out0(_handshake_buffer197_out0),
		.out0_valid(_handshake_buffer197_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer198(
		.in0(_handshake_cond_br21_outTrue),
		.in0_valid(_handshake_cond_br21_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork25_in0_ready),
		.in0_ready(_handshake_buffer198_in0_ready),
		.out0(_handshake_buffer198_out0),
		.out0_valid(_handshake_buffer198_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork24(
		.in0(_handshake_buffer197_out0),
		.in0_valid(_handshake_buffer197_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer200_in0_ready),
		.out1_ready(_handshake_buffer199_in0_ready),
		.in0_ready(_handshake_fork24_in0_ready),
		.out0(_handshake_fork24_out0),
		.out0_valid(_handshake_fork24_out0_valid),
		.out1(_handshake_fork24_out1),
		.out1_valid(_handshake_fork24_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer199(
		.in0(_handshake_fork24_out1),
		.in0_valid(_handshake_fork24_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli6_in0_ready),
		.in0_ready(_handshake_buffer199_in0_ready),
		.out0(_handshake_buffer199_out0),
		.out0_valid(_handshake_buffer199_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer200(
		.in0(_handshake_fork24_out0),
		.in0_valid(_handshake_fork24_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux11_in1_ready),
		.in0_ready(_handshake_buffer200_in0_ready),
		.out0(_handshake_buffer200_out0),
		.out0_valid(_handshake_buffer200_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork25(
		.in0(_handshake_buffer198_out0),
		.in0_valid(_handshake_buffer198_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer202_in0_ready),
		.out1_ready(_handshake_buffer201_in0_ready),
		.in0_ready(_handshake_fork25_in0_ready),
		.out0(_handshake_fork25_out0),
		.out0_valid(_handshake_fork25_out0_valid),
		.out1(_handshake_fork25_out1),
		.out1_valid(_handshake_fork25_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer201(
		.in0(_handshake_fork25_out1),
		.in0_valid(_handshake_fork25_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli2_in0_ready),
		.in0_ready(_handshake_buffer201_in0_ready),
		.out0(_handshake_buffer201_out0),
		.out0_valid(_handshake_buffer201_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer202(
		.in0(_handshake_fork25_out0),
		.in0_valid(_handshake_fork25_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux20_in1_ready),
		.in0_ready(_handshake_buffer202_in0_ready),
		.out0(_handshake_buffer202_out0),
		.out0_valid(_handshake_buffer202_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br22(
		.cond(_handshake_buffer175_out0),
		.cond_valid(_handshake_buffer175_out0_valid),
		.data(_handshake_buffer146_out0),
		.data_valid(_handshake_buffer146_out0_valid),
		.outTrue_ready(_handshake_buffer204_in0_ready),
		.outFalse_ready(_handshake_buffer203_in0_ready),
		.cond_ready(_handshake_cond_br22_cond_ready),
		.data_ready(_handshake_cond_br22_data_ready),
		.outTrue(_handshake_cond_br22_outTrue),
		.outTrue_valid(_handshake_cond_br22_outTrue_valid),
		.outFalse(_handshake_cond_br22_outFalse),
		.outFalse_valid(_handshake_cond_br22_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer203(
		.in0(_handshake_cond_br22_outFalse),
		.in0_valid(_handshake_cond_br22_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux12_in1_ready),
		.in0_ready(_handshake_buffer203_in0_ready),
		.out0(_handshake_buffer203_out0),
		.out0_valid(_handshake_buffer203_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer204(
		.in0(_handshake_cond_br22_outTrue),
		.in0_valid(_handshake_cond_br22_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux21_in1_ready),
		.in0_ready(_handshake_buffer204_in0_ready),
		.out0(_handshake_buffer204_out0),
		.out0_valid(_handshake_buffer204_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br23(
		.cond(_handshake_buffer176_out0),
		.cond_valid(_handshake_buffer176_out0_valid),
		.data(_handshake_buffer147_out0),
		.data_valid(_handshake_buffer147_out0_valid),
		.outTrue_ready(_handshake_buffer206_in0_ready),
		.outFalse_ready(_handshake_buffer205_in0_ready),
		.cond_ready(_handshake_cond_br23_cond_ready),
		.data_ready(_handshake_cond_br23_data_ready),
		.outTrue(_handshake_cond_br23_outTrue),
		.outTrue_valid(_handshake_cond_br23_outTrue_valid),
		.outFalse(_handshake_cond_br23_outFalse),
		.outFalse_valid(_handshake_cond_br23_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer205(
		.in0(_handshake_cond_br23_outFalse),
		.in0_valid(_handshake_cond_br23_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork26_in0_ready),
		.in0_ready(_handshake_buffer205_in0_ready),
		.out0(_handshake_buffer205_out0),
		.out0_valid(_handshake_buffer205_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer206(
		.in0(_handshake_cond_br23_outTrue),
		.in0_valid(_handshake_cond_br23_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux22_in1_ready),
		.in0_ready(_handshake_buffer206_in0_ready),
		.out0(_handshake_buffer206_out0),
		.out0_valid(_handshake_buffer206_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork26(
		.in0(_handshake_buffer205_out0),
		.in0_valid(_handshake_buffer205_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer208_in0_ready),
		.out1_ready(_handshake_buffer207_in0_ready),
		.in0_ready(_handshake_fork26_in0_ready),
		.out0(_handshake_fork26_out0),
		.out0_valid(_handshake_fork26_out0_valid),
		.out1(_handshake_fork26_out1),
		.out1_valid(_handshake_fork26_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer207(
		.in0(_handshake_fork26_out1),
		.in0_valid(_handshake_fork26_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi6_in1_ready),
		.in0_ready(_handshake_buffer207_in0_ready),
		.out0(_handshake_buffer207_out0),
		.out0_valid(_handshake_buffer207_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer208(
		.in0(_handshake_fork26_out0),
		.in0_valid(_handshake_fork26_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux13_in1_ready),
		.in0_ready(_handshake_buffer208_in0_ready),
		.out0(_handshake_buffer208_out0),
		.out0_valid(_handshake_buffer208_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br24(
		.cond(_handshake_buffer177_out0),
		.cond_valid(_handshake_buffer177_out0_valid),
		.data(_handshake_buffer148_out0),
		.data_valid(_handshake_buffer148_out0_valid),
		.outTrue_ready(_handshake_buffer210_in0_ready),
		.outFalse_ready(_handshake_buffer209_in0_ready),
		.cond_ready(_handshake_cond_br24_cond_ready),
		.data_ready(_handshake_cond_br24_data_ready),
		.outTrue(_handshake_cond_br24_outTrue),
		.outTrue_valid(_handshake_cond_br24_outTrue_valid),
		.outFalse(_handshake_cond_br24_outFalse),
		.outFalse_valid(_handshake_cond_br24_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer209(
		.in0(_handshake_cond_br24_outFalse),
		.in0_valid(_handshake_cond_br24_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork27_in0_ready),
		.in0_ready(_handshake_buffer209_in0_ready),
		.out0(_handshake_buffer209_out0),
		.out0_valid(_handshake_buffer209_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer210(
		.in0(_handshake_cond_br24_outTrue),
		.in0_valid(_handshake_cond_br24_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork28_in0_ready),
		.in0_ready(_handshake_buffer210_in0_ready),
		.out0(_handshake_buffer210_out0),
		.out0_valid(_handshake_buffer210_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork27(
		.in0(_handshake_buffer209_out0),
		.in0_valid(_handshake_buffer209_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer212_in0_ready),
		.out1_ready(_handshake_buffer211_in0_ready),
		.in0_ready(_handshake_fork27_in0_ready),
		.out0(_handshake_fork27_out0),
		.out0_valid(_handshake_fork27_out0_valid),
		.out1(_handshake_fork27_out1),
		.out1_valid(_handshake_fork27_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer211(
		.in0(_handshake_fork27_out1),
		.in0_valid(_handshake_fork27_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi6_in0_ready),
		.in0_ready(_handshake_buffer211_in0_ready),
		.out0(_handshake_buffer211_out0),
		.out0_valid(_handshake_buffer211_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer212(
		.in0(_handshake_fork27_out0),
		.in0_valid(_handshake_fork27_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi5_in1_ready),
		.in0_ready(_handshake_buffer212_in0_ready),
		.out0(_handshake_buffer212_out0),
		.out0_valid(_handshake_buffer212_out0_valid)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork28(
		.in0(_handshake_buffer210_out0),
		.in0_valid(_handshake_buffer210_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer214_in0_ready),
		.out1_ready(_handshake_buffer213_in0_ready),
		.in0_ready(_handshake_fork28_in0_ready),
		.out0(_handshake_fork28_out0),
		.out0_valid(_handshake_fork28_out0_valid),
		.out1(_handshake_fork28_out1),
		.out1_valid(_handshake_fork28_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer213(
		.in0(_handshake_fork28_out1),
		.in0_valid(_handshake_fork28_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi2_in1_ready),
		.in0_ready(_handshake_buffer213_in0_ready),
		.out0(_handshake_buffer213_out0),
		.out0_valid(_handshake_buffer213_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer214(
		.in0(_handshake_fork28_out0),
		.in0_valid(_handshake_fork28_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux23_in1_ready),
		.in0_ready(_handshake_buffer214_in0_ready),
		.out0(_handshake_buffer214_out0),
		.out0_valid(_handshake_buffer214_out0_valid)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br25(
		.cond(_handshake_buffer178_out0),
		.cond_valid(_handshake_buffer178_out0_valid),
		.data(_handshake_buffer151_out0),
		.data_valid(_handshake_buffer151_out0_valid),
		.outTrue_ready(_handshake_buffer215_in0_ready),
		.outFalse_ready(_handshake_sink9_in0_ready),
		.cond_ready(_handshake_cond_br25_cond_ready),
		.data_ready(_handshake_cond_br25_data_ready),
		.outTrue(_handshake_cond_br25_outTrue),
		.outTrue_valid(_handshake_cond_br25_outTrue_valid),
		.outFalse(_handshake_cond_br25_outFalse),
		.outFalse_valid(_handshake_cond_br25_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer215(
		.in0(_handshake_cond_br25_outTrue),
		.in0_valid(_handshake_cond_br25_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux24_in1_ready),
		.in0_ready(_handshake_buffer215_in0_ready),
		.out0(_handshake_buffer215_out0),
		.out0_valid(_handshake_buffer215_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink9(
		.in0(_handshake_cond_br25_outFalse),
		.in0_valid(_handshake_cond_br25_outFalse_valid),
		.in0_ready(_handshake_sink9_in0_ready)
	);
	handshake_cond_br_in_ui1_ui64_out_ui64_ui64 handshake_cond_br26(
		.cond(_handshake_buffer179_out0),
		.cond_valid(_handshake_buffer179_out0_valid),
		.data(_handshake_buffer152_out0),
		.data_valid(_handshake_buffer152_out0_valid),
		.outTrue_ready(_handshake_buffer216_in0_ready),
		.outFalse_ready(_handshake_sink10_in0_ready),
		.cond_ready(_handshake_cond_br26_cond_ready),
		.data_ready(_handshake_cond_br26_data_ready),
		.outTrue(_handshake_cond_br26_outTrue),
		.outTrue_valid(_handshake_cond_br26_outTrue_valid),
		.outFalse(_handshake_cond_br26_outFalse),
		.outFalse_valid(_handshake_cond_br26_outFalse_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer216(
		.in0(_handshake_cond_br26_outTrue),
		.in0_valid(_handshake_cond_br26_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork29_in0_ready),
		.in0_ready(_handshake_buffer216_in0_ready),
		.out0(_handshake_buffer216_out0),
		.out0_valid(_handshake_buffer216_out0_valid)
	);
	handshake_sink_in_ui64 handshake_sink10(
		.in0(_handshake_cond_br26_outFalse),
		.in0_valid(_handshake_cond_br26_outFalse_valid),
		.in0_ready(_handshake_sink10_in0_ready)
	);
	handshake_fork_in_ui64_out_ui64_ui64 handshake_fork29(
		.in0(_handshake_buffer216_out0),
		.in0_valid(_handshake_buffer216_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer218_in0_ready),
		.out1_ready(_handshake_buffer217_in0_ready),
		.in0_ready(_handshake_fork29_in0_ready),
		.out0(_handshake_fork29_out0),
		.out0_valid(_handshake_fork29_out0_valid),
		.out1(_handshake_fork29_out1),
		.out1_valid(_handshake_fork29_out1_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer217(
		.in0(_handshake_fork29_out1),
		.in0_valid(_handshake_fork29_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi4_in1_ready),
		.in0_ready(_handshake_buffer217_in0_ready),
		.out0(_handshake_buffer217_out0),
		.out0_valid(_handshake_buffer217_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer218(
		.in0(_handshake_fork29_out0),
		.in0_valid(_handshake_fork29_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux25_in1_ready),
		.in0_ready(_handshake_buffer218_in0_ready),
		.out0(_handshake_buffer218_out0),
		.out0_valid(_handshake_buffer218_out0_valid)
	);
	handshake_cond_br_in_ui1_2ins_2outs_ctrl handshake_cond_br27(
		.cond(_handshake_buffer180_out0),
		.cond_valid(_handshake_buffer180_out0_valid),
		.data_valid(_handshake_buffer154_out0_valid),
		.outTrue_ready(_handshake_buffer220_in0_ready),
		.outFalse_ready(_handshake_buffer219_in0_ready),
		.cond_ready(_handshake_cond_br27_cond_ready),
		.data_ready(_handshake_cond_br27_data_ready),
		.outTrue_valid(_handshake_cond_br27_outTrue_valid),
		.outFalse_valid(_handshake_cond_br27_outFalse_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer219(
		.in0_valid(_handshake_cond_br27_outFalse_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork30_in0_ready),
		.in0_ready(_handshake_buffer219_in0_ready),
		.out0_valid(_handshake_buffer219_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer220(
		.in0_valid(_handshake_cond_br27_outTrue_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_fork31_in0_ready),
		.in0_ready(_handshake_buffer220_in0_ready),
		.out0_valid(_handshake_buffer220_out0_valid)
	);
	handshake_fork_1ins_3outs_ctrl handshake_fork30(
		.in0_valid(_handshake_buffer219_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer223_in0_ready),
		.out1_ready(_handshake_buffer222_in0_ready),
		.out2_ready(_handshake_buffer221_in0_ready),
		.in0_ready(_handshake_fork30_in0_ready),
		.out0_valid(_handshake_fork30_out0_valid),
		.out1_valid(_handshake_fork30_out1_valid),
		.out2_valid(_handshake_fork30_out2_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer221(
		.in0_valid(_handshake_fork30_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant12_ctrl_ready),
		.in0_ready(_handshake_buffer221_in0_ready),
		.out0_valid(_handshake_buffer221_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer222(
		.in0_valid(_handshake_fork30_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join5_in0_ready),
		.in0_ready(_handshake_buffer222_in0_ready),
		.out0_valid(_handshake_buffer222_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer223(
		.in0_valid(_handshake_fork30_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_store0_ctrl_ready),
		.in0_ready(_handshake_buffer223_in0_ready),
		.out0_valid(_handshake_buffer223_out0_valid)
	);
	handshake_fork_1ins_5outs_ctrl handshake_fork31(
		.in0_valid(_handshake_buffer220_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_buffer228_in0_ready),
		.out1_ready(_handshake_buffer227_in0_ready),
		.out2_ready(_handshake_buffer226_in0_ready),
		.out3_ready(_handshake_buffer225_in0_ready),
		.out4_ready(_handshake_buffer224_in0_ready),
		.in0_ready(_handshake_fork31_in0_ready),
		.out0_valid(_handshake_fork31_out0_valid),
		.out1_valid(_handshake_fork31_out1_valid),
		.out2_valid(_handshake_fork31_out2_valid),
		.out3_valid(_handshake_fork31_out3_valid),
		.out4_valid(_handshake_fork31_out4_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer224(
		.in0_valid(_handshake_fork31_out4_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant10_ctrl_ready),
		.in0_ready(_handshake_buffer224_in0_ready),
		.out0_valid(_handshake_buffer224_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer225(
		.in0_valid(_handshake_fork31_out3_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_constant11_ctrl_ready),
		.in0_ready(_handshake_buffer225_in0_ready),
		.out0_valid(_handshake_buffer225_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer226(
		.in0_valid(_handshake_fork31_out2_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load1_ctrl_ready),
		.in0_ready(_handshake_buffer226_in0_ready),
		.out0_valid(_handshake_buffer226_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer227(
		.in0_valid(_handshake_fork31_out1_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_join4_in0_ready),
		.in0_ready(_handshake_buffer227_in0_ready),
		.out0_valid(_handshake_buffer227_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer228(
		.in0_valid(_handshake_fork31_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load2_ctrl_ready),
		.in0_ready(_handshake_buffer228_in0_ready),
		.out0_valid(_handshake_buffer228_out0_valid)
	);
	handshake_join_3ins_1outs_ctrl handshake_join4(
		.in0_valid(_handshake_buffer227_out0_valid),
		.in1_valid(_handshake_buffer23_out0_valid),
		.in2_valid(_handshake_buffer19_out0_valid),
		.out0_ready(_handshake_buffer229_in0_ready),
		.in0_ready(_handshake_join4_in0_ready),
		.in1_ready(_handshake_join4_in1_ready),
		.in2_ready(_handshake_join4_in2_ready),
		.out0_valid(_handshake_join4_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer229(
		.in0_valid(_handshake_join4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_control_merge1_in1_ready),
		.in0_ready(_handshake_buffer229_in0_ready),
		.out0_valid(_handshake_buffer229_out0_valid)
	);
	handshake_constant_c30_out_ui64 handshake_constant10(
		.ctrl_valid(_handshake_buffer224_out0_valid),
		.out0_ready(_handshake_buffer230_in0_ready),
		.ctrl_ready(_handshake_constant10_ctrl_ready),
		.out0(_handshake_constant10_out0),
		.out0_valid(_handshake_constant10_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer230(
		.in0(_handshake_constant10_out0),
		.in0_valid(_handshake_constant10_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli2_in1_ready),
		.in0_ready(_handshake_buffer230_in0_ready),
		.out0(_handshake_buffer230_out0),
		.out0_valid(_handshake_buffer230_out0_valid)
	);
	arith_muli_in_ui64_ui64_out_ui64 arith_muli2(
		.in0(_handshake_buffer201_out0),
		.in0_valid(_handshake_buffer201_out0_valid),
		.in1(_handshake_buffer230_out0),
		.in1_valid(_handshake_buffer230_out0_valid),
		.out0_ready(_handshake_buffer231_in0_ready),
		.in0_ready(_arith_muli2_in0_ready),
		.in1_ready(_arith_muli2_in1_ready),
		.out0(_arith_muli2_out0),
		.out0_valid(_arith_muli2_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer231(
		.in0(_arith_muli2_out0),
		.in0_valid(_arith_muli2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi1_in0_ready),
		.in0_ready(_handshake_buffer231_in0_ready),
		.out0(_handshake_buffer231_out0),
		.out0_valid(_handshake_buffer231_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi1(
		.in0(_handshake_buffer231_out0),
		.in0_valid(_handshake_buffer231_out0_valid),
		.in1(_handshake_buffer184_out0),
		.in1_valid(_handshake_buffer184_out0_valid),
		.out0_ready(_handshake_buffer232_in0_ready),
		.in0_ready(_arith_addi1_in0_ready),
		.in1_ready(_arith_addi1_in1_ready),
		.out0(_arith_addi1_out0),
		.out0_valid(_arith_addi1_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer232(
		.in0(_arith_addi1_out0),
		.in0_valid(_arith_addi1_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load1_addrIn0_ready),
		.in0_ready(_handshake_buffer232_in0_ready),
		.out0(_handshake_buffer232_out0),
		.out0_valid(_handshake_buffer232_out0_valid)
	);
	handshake_load_in_ui64_ui32_out_ui32_ui64 handshake_load1(
		.addrIn0(_handshake_buffer232_out0),
		.addrIn0_valid(_handshake_buffer232_out0_valid),
		.dataFromMem(_handshake_buffer22_out0),
		.dataFromMem_valid(_handshake_buffer22_out0_valid),
		.ctrl_valid(_handshake_buffer226_out0_valid),
		.dataOut_ready(_handshake_buffer234_in0_ready),
		.addrOut0_ready(_handshake_buffer233_in0_ready),
		.addrIn0_ready(_handshake_load1_addrIn0_ready),
		.dataFromMem_ready(_handshake_load1_dataFromMem_ready),
		.ctrl_ready(_handshake_load1_ctrl_ready),
		.dataOut(_handshake_load1_dataOut),
		.dataOut_valid(_handshake_load1_dataOut_valid),
		.addrOut0(_handshake_load1_addrOut0),
		.addrOut0_valid(_handshake_load1_addrOut0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer233(
		.in0(_handshake_load1_addrOut0),
		.in0_valid(_handshake_load1_addrOut0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_index_cast3_in0_ready),
		.in0_ready(_handshake_buffer233_in0_ready),
		.out0(_handshake_buffer233_out0),
		.out0_valid(_handshake_buffer233_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer234(
		.in0(_handshake_load1_dataOut),
		.in0_valid(_handshake_load1_dataOut_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli3_in1_ready),
		.in0_ready(_handshake_buffer234_in0_ready),
		.out0(_handshake_buffer234_out0),
		.out0_valid(_handshake_buffer234_out0_valid)
	);
	arith_muli_in_ui32_ui32_out_ui32 arith_muli3(
		.in0(_handshake_buffer189_out0),
		.in0_valid(_handshake_buffer189_out0_valid),
		.in1(_handshake_buffer234_out0),
		.in1_valid(_handshake_buffer234_out0_valid),
		.out0_ready(_handshake_buffer235_in0_ready),
		.in0_ready(_arith_muli3_in0_ready),
		.in1_ready(_arith_muli3_in1_ready),
		.out0(_arith_muli3_out0),
		.out0_valid(_arith_muli3_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer235(
		.in0(_arith_muli3_out0),
		.in0_valid(_arith_muli3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli5_in0_ready),
		.in0_ready(_handshake_buffer235_in0_ready),
		.out0(_handshake_buffer235_out0),
		.out0_valid(_handshake_buffer235_out0_valid)
	);
	handshake_constant_c30_out_ui64 handshake_constant11(
		.ctrl_valid(_handshake_buffer225_out0_valid),
		.out0_ready(_handshake_buffer236_in0_ready),
		.ctrl_ready(_handshake_constant11_ctrl_ready),
		.out0(_handshake_constant11_out0),
		.out0_valid(_handshake_constant11_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer236(
		.in0(_handshake_constant11_out0),
		.in0_valid(_handshake_constant11_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli4_in1_ready),
		.in0_ready(_handshake_buffer236_in0_ready),
		.out0(_handshake_buffer236_out0),
		.out0_valid(_handshake_buffer236_out0_valid)
	);
	arith_muli_in_ui64_ui64_out_ui64 arith_muli4(
		.in0(_handshake_buffer183_out0),
		.in0_valid(_handshake_buffer183_out0_valid),
		.in1(_handshake_buffer236_out0),
		.in1_valid(_handshake_buffer236_out0_valid),
		.out0_ready(_handshake_buffer237_in0_ready),
		.in0_ready(_arith_muli4_in0_ready),
		.in1_ready(_arith_muli4_in1_ready),
		.out0(_arith_muli4_out0),
		.out0_valid(_arith_muli4_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer237(
		.in0(_arith_muli4_out0),
		.in0_valid(_arith_muli4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi2_in0_ready),
		.in0_ready(_handshake_buffer237_in0_ready),
		.out0(_handshake_buffer237_out0),
		.out0_valid(_handshake_buffer237_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi2(
		.in0(_handshake_buffer237_out0),
		.in0_valid(_handshake_buffer237_out0_valid),
		.in1(_handshake_buffer213_out0),
		.in1_valid(_handshake_buffer213_out0_valid),
		.out0_ready(_handshake_buffer238_in0_ready),
		.in0_ready(_arith_addi2_in0_ready),
		.in1_ready(_arith_addi2_in1_ready),
		.out0(_arith_addi2_out0),
		.out0_valid(_arith_addi2_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer238(
		.in0(_arith_addi2_out0),
		.in0_valid(_arith_addi2_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_load2_addrIn0_ready),
		.in0_ready(_handshake_buffer238_in0_ready),
		.out0(_handshake_buffer238_out0),
		.out0_valid(_handshake_buffer238_out0_valid)
	);
	handshake_load_in_ui64_ui32_out_ui32_ui64 handshake_load2(
		.addrIn0(_handshake_buffer238_out0),
		.addrIn0_valid(_handshake_buffer238_out0_valid),
		.dataFromMem(_handshake_buffer18_out0),
		.dataFromMem_valid(_handshake_buffer18_out0_valid),
		.ctrl_valid(_handshake_buffer228_out0_valid),
		.dataOut_ready(_handshake_buffer240_in0_ready),
		.addrOut0_ready(_handshake_buffer239_in0_ready),
		.addrIn0_ready(_handshake_load2_addrIn0_ready),
		.dataFromMem_ready(_handshake_load2_dataFromMem_ready),
		.ctrl_ready(_handshake_load2_ctrl_ready),
		.dataOut(_handshake_load2_dataOut),
		.dataOut_valid(_handshake_load2_dataOut_valid),
		.addrOut0(_handshake_load2_addrOut0),
		.addrOut0_valid(_handshake_load2_addrOut0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer239(
		.in0(_handshake_load2_addrOut0),
		.in0_valid(_handshake_load2_addrOut0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_index_cast2_in0_ready),
		.in0_ready(_handshake_buffer239_in0_ready),
		.out0(_handshake_buffer239_out0),
		.out0_valid(_handshake_buffer239_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer240(
		.in0(_handshake_load2_dataOut),
		.in0_valid(_handshake_load2_dataOut_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli5_in1_ready),
		.in0_ready(_handshake_buffer240_in0_ready),
		.out0(_handshake_buffer240_out0),
		.out0_valid(_handshake_buffer240_out0_valid)
	);
	arith_muli_in_ui32_ui32_out_ui32 arith_muli5(
		.in0(_handshake_buffer235_out0),
		.in0_valid(_handshake_buffer235_out0_valid),
		.in1(_handshake_buffer240_out0),
		.in1_valid(_handshake_buffer240_out0_valid),
		.out0_ready(_handshake_buffer241_in0_ready),
		.in0_ready(_arith_muli5_in0_ready),
		.in1_ready(_arith_muli5_in1_ready),
		.out0(_arith_muli5_out0),
		.out0_valid(_arith_muli5_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer241(
		.in0(_arith_muli5_out0),
		.in0_valid(_arith_muli5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi3_in1_ready),
		.in0_ready(_handshake_buffer241_in0_ready),
		.out0(_handshake_buffer241_out0),
		.out0_valid(_handshake_buffer241_out0_valid)
	);
	arith_addi_in_ui32_ui32_out_ui32 arith_addi3(
		.in0(_handshake_buffer186_out0),
		.in0_valid(_handshake_buffer186_out0_valid),
		.in1(_handshake_buffer241_out0),
		.in1_valid(_handshake_buffer241_out0_valid),
		.out0_ready(_handshake_buffer242_in0_ready),
		.in0_ready(_arith_addi3_in0_ready),
		.in1_ready(_arith_addi3_in1_ready),
		.out0(_arith_addi3_out0),
		.out0_valid(_arith_addi3_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer242(
		.in0(_arith_addi3_out0),
		.in0_valid(_arith_addi3_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux15_in1_ready),
		.in0_ready(_handshake_buffer242_in0_ready),
		.out0(_handshake_buffer242_out0),
		.out0_valid(_handshake_buffer242_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi4(
		.in0(_handshake_buffer182_out0),
		.in0_valid(_handshake_buffer182_out0_valid),
		.in1(_handshake_buffer217_out0),
		.in1_valid(_handshake_buffer217_out0_valid),
		.out0_ready(_handshake_buffer243_in0_ready),
		.in0_ready(_arith_addi4_in0_ready),
		.in1_ready(_arith_addi4_in1_ready),
		.out0(_arith_addi4_out0),
		.out0_valid(_arith_addi4_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer243(
		.in0(_arith_addi4_out0),
		.in0_valid(_arith_addi4_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux14_in1_ready),
		.in0_ready(_handshake_buffer243_in0_ready),
		.out0(_handshake_buffer243_out0),
		.out0_valid(_handshake_buffer243_out0_valid)
	);
	handshake_join_2ins_1outs_ctrl handshake_join5(
		.in0_valid(_handshake_buffer222_out0_valid),
		.in1_valid(_handshake_buffer1_out0_valid),
		.out0_ready(_handshake_buffer244_in0_ready),
		.in0_ready(_handshake_join5_in0_ready),
		.in1_ready(_handshake_join5_in1_ready),
		.out0_valid(_handshake_join5_out0_valid)
	);
	handshake_buffer_2slots_seq_1ins_1outs_ctrl handshake_buffer244(
		.in0_valid(_handshake_join5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_control_merge0_in1_ready),
		.in0_ready(_handshake_buffer244_in0_ready),
		.out0_valid(_handshake_buffer244_out0_valid)
	);
	handshake_constant_c30_out_ui64 handshake_constant12(
		.ctrl_valid(_handshake_buffer221_out0_valid),
		.out0_ready(_handshake_buffer245_in0_ready),
		.ctrl_ready(_handshake_constant12_ctrl_ready),
		.out0(_handshake_constant12_out0),
		.out0_valid(_handshake_constant12_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer245(
		.in0(_handshake_constant12_out0),
		.in0_valid(_handshake_constant12_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_muli6_in1_ready),
		.in0_ready(_handshake_buffer245_in0_ready),
		.out0(_handshake_buffer245_out0),
		.out0_valid(_handshake_buffer245_out0_valid)
	);
	arith_muli_in_ui64_ui64_out_ui64 arith_muli6(
		.in0(_handshake_buffer199_out0),
		.in0_valid(_handshake_buffer199_out0_valid),
		.in1(_handshake_buffer245_out0),
		.in1_valid(_handshake_buffer245_out0_valid),
		.out0_ready(_handshake_buffer246_in0_ready),
		.in0_ready(_arith_muli6_in0_ready),
		.in1_ready(_arith_muli6_in1_ready),
		.out0(_arith_muli6_out0),
		.out0_valid(_arith_muli6_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer246(
		.in0(_arith_muli6_out0),
		.in0_valid(_arith_muli6_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_addi5_in0_ready),
		.in0_ready(_handshake_buffer246_in0_ready),
		.out0(_handshake_buffer246_out0),
		.out0_valid(_handshake_buffer246_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi5(
		.in0(_handshake_buffer246_out0),
		.in0_valid(_handshake_buffer246_out0_valid),
		.in1(_handshake_buffer212_out0),
		.in1_valid(_handshake_buffer212_out0_valid),
		.out0_ready(_handshake_buffer247_in0_ready),
		.in0_ready(_arith_addi5_in0_ready),
		.in1_ready(_arith_addi5_in1_ready),
		.out0(_arith_addi5_out0),
		.out0_valid(_arith_addi5_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer247(
		.in0(_arith_addi5_out0),
		.in0_valid(_arith_addi5_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_store0_addrIn0_ready),
		.in0_ready(_handshake_buffer247_in0_ready),
		.out0(_handshake_buffer247_out0),
		.out0_valid(_handshake_buffer247_out0_valid)
	);
	handshake_store_in_ui64_ui32_out_ui32_ui64 handshake_store0(
		.addrIn0(_handshake_buffer247_out0),
		.addrIn0_valid(_handshake_buffer247_out0_valid),
		.dataIn(_handshake_buffer185_out0),
		.dataIn_valid(_handshake_buffer185_out0_valid),
		.ctrl_valid(_handshake_buffer223_out0_valid),
		.dataToMem_ready(_handshake_buffer249_in0_ready),
		.addrOut0_ready(_handshake_buffer248_in0_ready),
		.addrIn0_ready(_handshake_store0_addrIn0_ready),
		.dataIn_ready(_handshake_store0_dataIn_ready),
		.ctrl_ready(_handshake_store0_ctrl_ready),
		.dataToMem(_handshake_store0_dataToMem),
		.dataToMem_valid(_handshake_store0_dataToMem_valid),
		.addrOut0(_handshake_store0_addrOut0),
		.addrOut0_valid(_handshake_store0_addrOut0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer248(
		.in0(_handshake_store0_addrOut0),
		.in0_valid(_handshake_store0_addrOut0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_arith_index_cast1_in0_ready),
		.in0_ready(_handshake_buffer248_in0_ready),
		.out0(_handshake_buffer248_out0),
		.out0_valid(_handshake_buffer248_out0_valid)
	);
	handshake_buffer_in_ui32_out_ui32_2slots_seq handshake_buffer249(
		.in0(_handshake_store0_dataToMem),
		.in0_valid(_handshake_store0_dataToMem_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_hw_struct_create0_in1_ready),
		.in0_ready(_handshake_buffer249_in0_ready),
		.out0(_handshake_buffer249_out0),
		.out0_valid(_handshake_buffer249_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi6(
		.in0(_handshake_buffer211_out0),
		.in0_valid(_handshake_buffer211_out0_valid),
		.in1(_handshake_buffer207_out0),
		.in1_valid(_handshake_buffer207_out0_valid),
		.out0_ready(_handshake_buffer250_in0_ready),
		.in0_ready(_arith_addi6_in0_ready),
		.in1_ready(_arith_addi6_in1_ready),
		.out0(_arith_addi6_out0),
		.out0_valid(_arith_addi6_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer250(
		.in0(_arith_addi6_out0),
		.in0_valid(_arith_addi6_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux6_in1_ready),
		.in0_ready(_handshake_buffer250_in0_ready),
		.out0(_handshake_buffer250_out0),
		.out0_valid(_handshake_buffer250_out0_valid)
	);
	arith_addi_in_ui64_ui64_out_ui64 arith_addi7(
		.in0(_handshake_buffer113_out0),
		.in0_valid(_handshake_buffer113_out0_valid),
		.in1(_handshake_buffer111_out0),
		.in1_valid(_handshake_buffer111_out0_valid),
		.out0_ready(_handshake_buffer251_in0_ready),
		.in0_ready(_arith_addi7_in0_ready),
		.in1_ready(_arith_addi7_in1_ready),
		.out0(_arith_addi7_out0),
		.out0_valid(_arith_addi7_out0_valid)
	);
	handshake_buffer_in_ui64_out_ui64_2slots_seq handshake_buffer251(
		.in0(_arith_addi7_out0),
		.in0_valid(_arith_addi7_out0_valid),
		.clock(clock),
		.reset(reset),
		.out0_ready(_handshake_mux1_in1_ready),
		.in0_ready(_handshake_buffer251_in0_ready),
		.out0(_handshake_buffer251_out0),
		.out0_valid(_handshake_buffer251_out0_valid)
	);
endmodule
