module LUT4AB_switch_matrix #(
    parameter NoConfigBits = 1329
)(
    output N2BEGb0,
    output N2BEGb1,
    output N2BEGb2,
    output N2BEGb3,
    output N2BEGb4,
    output N2BEGb5,
    output N2BEGb6,
    output N2BEGb7,
    output E2BEGb0,
    output E2BEGb1,
    output E2BEGb2,
    output E2BEGb3,
    output E2BEGb4,
    output E2BEGb5,
    output E2BEGb6,
    output E2BEGb7,
    output S2BEGb0,
    output S2BEGb1,
    output S2BEGb2,
    output S2BEGb3,
    output S2BEGb4,
    output S2BEGb5,
    output S2BEGb6,
    output S2BEGb7,
    output W2BEGb0,
    output W2BEGb1,
    output W2BEGb2,
    output W2BEGb3,
    output W2BEGb4,
    output W2BEGb5,
    output W2BEGb6,
    output W2BEGb7,
    output J2MID_ABa_BEG0,
    output J2MID_ABa_BEG1,
    output J2MID_ABa_BEG2,
    output J2MID_ABa_BEG3,
    output J2MID_CDa_BEG0,
    output J2MID_CDa_BEG1,
    output J2MID_CDa_BEG2,
    output J2MID_CDa_BEG3,
    output J2MID_EFa_BEG0,
    output J2MID_EFa_BEG1,
    output J2MID_EFa_BEG2,
    output J2MID_EFa_BEG3,
    output J2MID_GHa_BEG0,
    output J2MID_GHa_BEG1,
    output J2MID_GHa_BEG2,
    output J2MID_GHa_BEG3,
    output J2MID_ABb_BEG0,
    output J2MID_ABb_BEG1,
    output J2MID_ABb_BEG2,
    output J2MID_ABb_BEG3,
    output J2MID_CDb_BEG0,
    output J2MID_CDb_BEG1,
    output J2MID_CDb_BEG2,
    output J2MID_CDb_BEG3,
    output J2MID_EFb_BEG0,
    output J2MID_EFb_BEG1,
    output J2MID_EFb_BEG2,
    output J2MID_EFb_BEG3,
    output J2MID_GHb_BEG0,
    output J2MID_GHb_BEG1,
    output J2MID_GHb_BEG2,
    output J2MID_GHb_BEG3,
    output J2END_AB_BEG0,
    output J2END_AB_BEG1,
    output J2END_AB_BEG2,
    output J2END_AB_BEG3,
    output J2END_CD_BEG0,
    output J2END_CD_BEG1,
    output J2END_CD_BEG2,
    output J2END_CD_BEG3,
    output J2END_EF_BEG0,
    output J2END_EF_BEG1,
    output J2END_EF_BEG2,
    output J2END_EF_BEG3,
    output J2END_GH_BEG0,
    output J2END_GH_BEG1,
    output J2END_GH_BEG2,
    output J2END_GH_BEG3,
    output J_l_AB_BEG0,
    output J_l_AB_BEG1,
    output J_l_AB_BEG2,
    output J_l_AB_BEG3,
    output J_l_CD_BEG0,
    output J_l_CD_BEG1,
    output J_l_CD_BEG2,
    output J_l_CD_BEG3,
    output J_l_EF_BEG0,
    output J_l_EF_BEG1,
    output J_l_EF_BEG2,
    output J_l_EF_BEG3,
    output J_l_GH_BEG0,
    output J_l_GH_BEG1,
    output J_l_GH_BEG2,
    output J_l_GH_BEG3,
    output LA_I0,
    output LB_I0,
    output LA_I1,
    output LB_I1,
    output LA_I2,
    output LB_I2,
    output LA_I3,
    output LB_I3,
    output LC_I0,
    output LD_I0,
    output LC_I1,
    output LD_I1,
    output LC_I2,
    output LD_I2,
    output LC_I3,
    output LD_I3,
    output LE_I0,
    output LF_I0,
    output LE_I1,
    output LF_I1,
    output LE_I2,
    output LF_I2,
    output LE_I3,
    output LF_I3,
    output LG_I0,
    output LH_I0,
    output LG_I1,
    output LH_I1,
    output LG_I2,
    output LH_I2,
    output LG_I3,
    output LH_I3,
    output JN2BEG0,
    output JN2BEG1,
    output JN2BEG2,
    output JN2BEG3,
    output JN2BEG4,
    output JN2BEG5,
    output JN2BEG6,
    output JN2BEG7,
    output JE2BEG0,
    output JE2BEG1,
    output JE2BEG2,
    output JE2BEG3,
    output JE2BEG4,
    output JE2BEG5,
    output JE2BEG6,
    output JE2BEG7,
    output JS2BEG0,
    output JS2BEG1,
    output JS2BEG2,
    output JS2BEG3,
    output JS2BEG4,
    output JS2BEG5,
    output JS2BEG6,
    output JS2BEG7,
    output JW2BEG0,
    output JW2BEG1,
    output JW2BEG2,
    output JW2BEG3,
    output JW2BEG4,
    output JW2BEG5,
    output JW2BEG6,
    output JW2BEG7,
    output N2BEG0,
    output N2BEG1,
    output N2BEG2,
    output N2BEG3,
    output N2BEG4,
    output N2BEG5,
    output N2BEG6,
    output N2BEG7,
    output E2BEG0,
    output E2BEG1,
    output E2BEG2,
    output E2BEG3,
    output E2BEG4,
    output E2BEG5,
    output E2BEG6,
    output E2BEG7,
    output S2BEG0,
    output S2BEG1,
    output S2BEG2,
    output S2BEG3,
    output S2BEG4,
    output S2BEG5,
    output S2BEG6,
    output S2BEG7,
    output W2BEG1,
    output W2BEG2,
    output W2BEG5,
    output W2BEG6,
    output W2BEG0,
    output W2BEG3,
    output W2BEG4,
    output W2BEG7,
    output N1BEG0,
    output N1BEG1,
    output N1BEG2,
    output N1BEG3,
    output E1BEG0,
    output E1BEG1,
    output E1BEG2,
    output E1BEG3,
    output S1BEG0,
    output S1BEG1,
    output S1BEG2,
    output S1BEG3,
    output W1BEG0,
    output W1BEG1,
    output W1BEG2,
    output W1BEG3,
    output N4BEG0,
    output N4BEG1,
    output N4BEG2,
    output N4BEG3,
    output S4BEG0,
    output S4BEG1,
    output S4BEG2,
    output S4BEG3,
    output E6BEG0,
    output E6BEG1,
    output W6BEG0,
    output W6BEG1,
    output EE4BEG0,
    output EE4BEG1,
    output EE4BEG2,
    output EE4BEG3,
    output WW4BEG0,
    output WW4BEG1,
    output WW4BEG2,
    output WW4BEG3,
    output NN4BEG0,
    output NN4BEG1,
    output NN4BEG2,
    output NN4BEG3,
    output SS4BEG0,
    output SS4BEG1,
    output SS4BEG2,
    output SS4BEG3,
    output A,
    output B,
    output C,
    output D,
    output E,
    output F,
    output G,
    output H,
    output S0,
    output S1,
    output S2,
    output S3,
    output LA_Ci,
    output LB_Ci,
    output LC_Ci,
    output LD_Ci,
    output LE_Ci,
    output LF_Ci,
    output LG_Ci,
    output LH_Ci,
    output Co0,
    output J_SR_BEG0,
    output J_EN_BEG0,
    output LA_SR,
    output LB_SR,
    output LC_SR,
    output LD_SR,
    output LE_SR,
    output LF_SR,
    output LG_SR,
    output LH_SR,
    output LA_EN,
    output LB_EN,
    output LC_EN,
    output LD_EN,
    output LE_EN,
    output LF_EN,
    output LG_EN,
    output LH_EN,
    input N2MID0,
    input N2MID1,
    input N2MID2,
    input N2MID3,
    input N2MID4,
    input N2MID5,
    input N2MID6,
    input N2MID7,
    input E2MID0,
    input E2MID1,
    input E2MID2,
    input E2MID3,
    input E2MID4,
    input E2MID5,
    input E2MID6,
    input E2MID7,
    input S2MID0,
    input S2MID1,
    input S2MID2,
    input S2MID3,
    input S2MID4,
    input S2MID5,
    input S2MID6,
    input S2MID7,
    input W2MID0,
    input W2MID1,
    input W2MID2,
    input W2MID3,
    input W2MID4,
    input W2MID5,
    input W2MID6,
    input W2MID7,
    input JN2END3,
    input JE2END3,
    input JS2END3,
    input JW2END3,
    input JN2END4,
    input JE2END4,
    input JS2END4,
    input JW2END4,
    input JN2END5,
    input JE2END5,
    input JS2END5,
    input JW2END5,
    input JN2END6,
    input JE2END6,
    input JS2END6,
    input JW2END6,
    input E2END6,
    input N2END6,
    input SS4END3,
    input W2END6,
    input E2END2,
    input NN4END0,
    input S2END2,
    input W2END2,
    input EE4END0,
    input N2END4,
    input S2END4,
    input W2END4,
    input E2END0,
    input N2END0,
    input S2END0,
    input WW4END3,
    input NN4END3,
    input S2END6,
    input N2END2,
    input WW4END2,
    input E2END4,
    input SS4END2,
    input EE4END1,
    input W2END0,
    input EE4END2,
    input N2END7,
    input S2END7,
    input W2END7,
    input E2END3,
    input N2END3,
    input S2END3,
    input WW4END1,
    input E2END5,
    input N2END5,
    input SS4END1,
    input W2END5,
    input E2END1,
    input NN4END2,
    input S2END1,
    input W2END1,
    input E2END7,
    input WW4END0,
    input SS4END0,
    input W2END3,
    input NN4END1,
    input S2END5,
    input EE4END3,
    input N2END1,
    input JN2END1,
    input S4END3,
    input JE2END1,
    input S4END2,
    input E6END1,
    input N4END1,
    input JS2END1,
    input W6END1,
    input E6END0,
    input N4END0,
    input S4END0,
    input JW2END1,
    input JN2END2,
    input N4END2,
    input JE2END2,
    input S4END1,
    input JS2END2,
    input JW2END2,
    input W6END0,
    input N4END3,
    input J2MID_ABa_END0,
    input J2MID_ABb_END0,
    input J2END_AB_END0,
    input J_l_AB_END0,
    input J2MID_ABa_END1,
    input J2MID_ABb_END1,
    input J2END_AB_END1,
    input J_l_AB_END1,
    input J2MID_ABa_END2,
    input J2MID_ABb_END2,
    input J2END_AB_END2,
    input J_l_AB_END2,
    input J2MID_ABa_END3,
    input J2MID_ABb_END3,
    input J2END_AB_END3,
    input J_l_AB_END3,
    input J2MID_CDa_END0,
    input J2MID_CDb_END0,
    input J2END_CD_END0,
    input J_l_CD_END0,
    input J2MID_CDa_END1,
    input J2MID_CDb_END1,
    input J2END_CD_END1,
    input J_l_CD_END1,
    input J2MID_CDa_END2,
    input J2MID_CDb_END2,
    input J2END_CD_END2,
    input J_l_CD_END2,
    input J2MID_CDa_END3,
    input J2MID_CDb_END3,
    input J2END_CD_END3,
    input J_l_CD_END3,
    input J2MID_EFa_END0,
    input J2MID_EFb_END0,
    input J2END_EF_END0,
    input J_l_EF_END0,
    input J2MID_EFa_END1,
    input J2MID_EFb_END1,
    input J2END_EF_END1,
    input J_l_EF_END1,
    input J2MID_EFa_END2,
    input J2MID_EFb_END2,
    input J2END_EF_END2,
    input J_l_EF_END2,
    input J2MID_EFa_END3,
    input J2MID_EFb_END3,
    input J2END_EF_END3,
    input J_l_EF_END3,
    input J2MID_GHa_END0,
    input J2MID_GHb_END0,
    input J2END_GH_END0,
    input J_l_GH_END0,
    input J2MID_GHa_END1,
    input J2MID_GHb_END1,
    input J2END_GH_END1,
    input J_l_GH_END1,
    input J2MID_GHa_END2,
    input J2MID_GHb_END2,
    input J2END_GH_END2,
    input J_l_GH_END2,
    input J2MID_GHa_END3,
    input J2MID_GHb_END3,
    input J2END_GH_END3,
    input J_l_GH_END3,
    input E1END3,
    input LB_O,
    input LC_O,
    input LD_O,
    input LE_O,
    input LF_O,
    input LG_O,
    input LH_O,
    input M_AB,
    input LA_O,
    input E1END0,
    input M_AD,
    input E1END1,
    input M_AH,
    input E1END2,
    input M_EF,
    input W1END3,
    input N1END1,
    input S1END1,
    input W1END1,
    input W1END0,
    input N1END2,
    input S1END2,
    input W1END2,
    input N1END3,
    input S1END3,
    input N1END0,
    input S1END0,
    input JN2END0,
    input JN2END7,
    input JE2END0,
    input JE2END7,
    input JS2END0,
    input JS2END7,
    input JW2END0,
    input JW2END7,
    input Ci0,
    input LA_Co,
    input LB_Co,
    input LC_Co,
    input LD_Co,
    input LE_Co,
    input LF_Co,
    input LG_Co,
    input LH_Co,
    input J_SR_END0,
    input GND0,
    input J_EN_END0,
    input VCC0,
    input [NoConfigBits - 1:0] ConfigBits,
    input [NoConfigBits - 1:0] ConfigBits_N
);

localparam reg GND0 = 0;localparam reg GND = 0;localparam reg VCC0 = 1;localparam reg VCC = 1;localparam reg VDD0 = 1;localparam reg VDD = 1;// switch matrix multiplexer N2BEGb0 MUX-1assign N2BEGb0 = N2MID0;// switch matrix multiplexer N2BEGb1 MUX-1assign N2BEGb1 = N2MID1;// switch matrix multiplexer N2BEGb2 MUX-1assign N2BEGb2 = N2MID2;// switch matrix multiplexer N2BEGb3 MUX-1assign N2BEGb3 = N2MID3;// switch matrix multiplexer N2BEGb4 MUX-1assign N2BEGb4 = N2MID4;// switch matrix multiplexer N2BEGb5 MUX-1assign N2BEGb5 = N2MID5;// switch matrix multiplexer N2BEGb6 MUX-1assign N2BEGb6 = N2MID6;// switch matrix multiplexer N2BEGb7 MUX-1assign N2BEGb7 = N2MID7;// switch matrix multiplexer E2BEGb0 MUX-1assign E2BEGb0 = E2MID0;// switch matrix multiplexer E2BEGb1 MUX-1assign E2BEGb1 = E2MID1;// switch matrix multiplexer E2BEGb2 MUX-1assign E2BEGb2 = E2MID2;// switch matrix multiplexer E2BEGb3 MUX-1assign E2BEGb3 = E2MID3;// switch matrix multiplexer E2BEGb4 MUX-1assign E2BEGb4 = E2MID4;// switch matrix multiplexer E2BEGb5 MUX-1assign E2BEGb5 = E2MID5;// switch matrix multiplexer E2BEGb6 MUX-1assign E2BEGb6 = E2MID6;// switch matrix multiplexer E2BEGb7 MUX-1assign E2BEGb7 = E2MID7;// switch matrix multiplexer S2BEGb0 MUX-1assign S2BEGb0 = S2MID0;// switch matrix multiplexer S2BEGb1 MUX-1assign S2BEGb1 = S2MID1;// switch matrix multiplexer S2BEGb2 MUX-1assign S2BEGb2 = S2MID2;// switch matrix multiplexer S2BEGb3 MUX-1assign S2BEGb3 = S2MID3;// switch matrix multiplexer S2BEGb4 MUX-1assign S2BEGb4 = S2MID4;// switch matrix multiplexer S2BEGb5 MUX-1assign S2BEGb5 = S2MID5;// switch matrix multiplexer S2BEGb6 MUX-1assign S2BEGb6 = S2MID6;// switch matrix multiplexer S2BEGb7 MUX-1assign S2BEGb7 = S2MID7;// switch matrix multiplexer W2BEGb0 MUX-1assign W2BEGb0 = W2MID0;// switch matrix multiplexer W2BEGb1 MUX-1assign W2BEGb1 = W2MID1;// switch matrix multiplexer W2BEGb2 MUX-1assign W2BEGb2 = W2MID2;// switch matrix multiplexer W2BEGb3 MUX-1assign W2BEGb3 = W2MID3;// switch matrix multiplexer W2BEGb4 MUX-1assign W2BEGb4 = W2MID4;// switch matrix multiplexer W2BEGb5 MUX-1assign W2BEGb5 = W2MID5;// switch matrix multiplexer W2BEGb6 MUX-1assign W2BEGb6 = W2MID6;// switch matrix multiplexer W2BEGb7 MUX-1assign W2BEGb7 = W2MID7;// switch matrix multiplexer J2MID_ABa_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABa_BEG0 (
    .A0(W2MID6),
    .A1(S2MID6),
    .A2(N2MID6),
    .A3(JN2END3),
    .S0(ConfigBits[0]),
    .S0N(ConfigBits_N[0]),
    .S1(ConfigBits[1]),
    .S1N(ConfigBits_N[1]),
    .X(J2MID_ABa_BEG0)
);
// switch matrix multiplexer J2MID_ABa_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABa_BEG1 (
    .A0(W2MID2),
    .A1(S2MID2),
    .A2(JE2END3),
    .A3(E2MID2),
    .S0(ConfigBits[2]),
    .S0N(ConfigBits_N[2]),
    .S1(ConfigBits[3]),
    .S1N(ConfigBits_N[3]),
    .X(J2MID_ABa_BEG1)
);
// switch matrix multiplexer J2MID_ABa_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABa_BEG2 (
    .A0(W2MID4),
    .A1(JS2END3),
    .A2(N2MID4),
    .A3(E2MID4),
    .S0(ConfigBits[4]),
    .S0N(ConfigBits_N[4]),
    .S1(ConfigBits[5]),
    .S1N(ConfigBits_N[5]),
    .X(J2MID_ABa_BEG2)
);
// switch matrix multiplexer J2MID_ABa_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABa_BEG3 (
    .A0(JW2END3),
    .A1(S2MID0),
    .A2(N2MID0),
    .A3(E2MID0),
    .S0(ConfigBits[6]),
    .S0N(ConfigBits_N[6]),
    .S1(ConfigBits[7]),
    .S1N(ConfigBits_N[7]),
    .X(J2MID_ABa_BEG3)
);
// switch matrix multiplexer J2MID_CDa_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDa_BEG0 (
    .A0(W2MID6),
    .A1(S2MID6),
    .A2(JN2END4),
    .A3(E2MID6),
    .S0(ConfigBits[8]),
    .S0N(ConfigBits_N[8]),
    .S1(ConfigBits[9]),
    .S1N(ConfigBits_N[9]),
    .X(J2MID_CDa_BEG0)
);
// switch matrix multiplexer J2MID_CDa_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDa_BEG1 (
    .A0(W2MID2),
    .A1(JE2END4),
    .A2(N2MID2),
    .A3(E2MID2),
    .S0(ConfigBits[10]),
    .S0N(ConfigBits_N[10]),
    .S1(ConfigBits[11]),
    .S1N(ConfigBits_N[11]),
    .X(J2MID_CDa_BEG1)
);
// switch matrix multiplexer J2MID_CDa_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDa_BEG2 (
    .A0(JS2END4),
    .A1(S2MID4),
    .A2(N2MID4),
    .A3(E2MID4),
    .S0(ConfigBits[12]),
    .S0N(ConfigBits_N[12]),
    .S1(ConfigBits[13]),
    .S1N(ConfigBits_N[13]),
    .X(J2MID_CDa_BEG2)
);
// switch matrix multiplexer J2MID_CDa_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDa_BEG3 (
    .A0(W2MID0),
    .A1(S2MID0),
    .A2(N2MID0),
    .A3(JW2END4),
    .S0(ConfigBits[14]),
    .S0N(ConfigBits_N[14]),
    .S1(ConfigBits[15]),
    .S1N(ConfigBits_N[15]),
    .X(J2MID_CDa_BEG3)
);
// switch matrix multiplexer J2MID_EFa_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFa_BEG0 (
    .A0(W2MID6),
    .A1(JN2END5),
    .A2(N2MID6),
    .A3(E2MID6),
    .S0(ConfigBits[16]),
    .S0N(ConfigBits_N[16]),
    .S1(ConfigBits[17]),
    .S1N(ConfigBits_N[17]),
    .X(J2MID_EFa_BEG0)
);
// switch matrix multiplexer J2MID_EFa_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFa_BEG1 (
    .A0(JE2END5),
    .A1(S2MID2),
    .A2(N2MID2),
    .A3(E2MID2),
    .S0(ConfigBits[18]),
    .S0N(ConfigBits_N[18]),
    .S1(ConfigBits[19]),
    .S1N(ConfigBits_N[19]),
    .X(J2MID_EFa_BEG1)
);
// switch matrix multiplexer J2MID_EFa_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFa_BEG2 (
    .A0(W2MID4),
    .A1(S2MID4),
    .A2(N2MID4),
    .A3(JS2END5),
    .S0(ConfigBits[20]),
    .S0N(ConfigBits_N[20]),
    .S1(ConfigBits[21]),
    .S1N(ConfigBits_N[21]),
    .X(J2MID_EFa_BEG2)
);
// switch matrix multiplexer J2MID_EFa_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFa_BEG3 (
    .A0(W2MID0),
    .A1(S2MID0),
    .A2(JW2END5),
    .A3(E2MID0),
    .S0(ConfigBits[22]),
    .S0N(ConfigBits_N[22]),
    .S1(ConfigBits[23]),
    .S1N(ConfigBits_N[23]),
    .X(J2MID_EFa_BEG3)
);
// switch matrix multiplexer J2MID_GHa_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHa_BEG0 (
    .A0(JN2END6),
    .A1(S2MID6),
    .A2(N2MID6),
    .A3(E2MID6),
    .S0(ConfigBits[24]),
    .S0N(ConfigBits_N[24]),
    .S1(ConfigBits[25]),
    .S1N(ConfigBits_N[25]),
    .X(J2MID_GHa_BEG0)
);
// switch matrix multiplexer J2MID_GHa_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHa_BEG1 (
    .A0(W2MID2),
    .A1(S2MID2),
    .A2(N2MID2),
    .A3(JE2END6),
    .S0(ConfigBits[26]),
    .S0N(ConfigBits_N[26]),
    .S1(ConfigBits[27]),
    .S1N(ConfigBits_N[27]),
    .X(J2MID_GHa_BEG1)
);
// switch matrix multiplexer J2MID_GHa_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHa_BEG2 (
    .A0(W2MID4),
    .A1(S2MID4),
    .A2(JS2END6),
    .A3(E2MID4),
    .S0(ConfigBits[28]),
    .S0N(ConfigBits_N[28]),
    .S1(ConfigBits[29]),
    .S1N(ConfigBits_N[29]),
    .X(J2MID_GHa_BEG2)
);
// switch matrix multiplexer J2MID_GHa_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHa_BEG3 (
    .A0(W2MID0),
    .A1(JW2END6),
    .A2(N2MID0),
    .A3(E2MID0),
    .S0(ConfigBits[30]),
    .S0N(ConfigBits_N[30]),
    .S1(ConfigBits[31]),
    .S1N(ConfigBits_N[31]),
    .X(J2MID_GHa_BEG3)
);
// switch matrix multiplexer J2MID_ABb_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABb_BEG0 (
    .A0(W2MID7),
    .A1(S2MID7),
    .A2(N2MID7),
    .A3(E2MID7),
    .S0(ConfigBits[32]),
    .S0N(ConfigBits_N[32]),
    .S1(ConfigBits[33]),
    .S1N(ConfigBits_N[33]),
    .X(J2MID_ABb_BEG0)
);
// switch matrix multiplexer J2MID_ABb_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABb_BEG1 (
    .A0(W2MID3),
    .A1(S2MID3),
    .A2(N2MID3),
    .A3(E2MID3),
    .S0(ConfigBits[34]),
    .S0N(ConfigBits_N[34]),
    .S1(ConfigBits[35]),
    .S1N(ConfigBits_N[35]),
    .X(J2MID_ABb_BEG1)
);
// switch matrix multiplexer J2MID_ABb_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABb_BEG2 (
    .A0(W2MID5),
    .A1(S2MID5),
    .A2(N2MID5),
    .A3(E2MID5),
    .S0(ConfigBits[36]),
    .S0N(ConfigBits_N[36]),
    .S1(ConfigBits[37]),
    .S1N(ConfigBits_N[37]),
    .X(J2MID_ABb_BEG2)
);
// switch matrix multiplexer J2MID_ABb_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_ABb_BEG3 (
    .A0(W2MID1),
    .A1(S2MID1),
    .A2(N2MID1),
    .A3(E2MID1),
    .S0(ConfigBits[38]),
    .S0N(ConfigBits_N[38]),
    .S1(ConfigBits[39]),
    .S1N(ConfigBits_N[39]),
    .X(J2MID_ABb_BEG3)
);
// switch matrix multiplexer J2MID_CDb_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDb_BEG0 (
    .A0(W2MID7),
    .A1(S2MID7),
    .A2(N2MID7),
    .A3(E2MID7),
    .S0(ConfigBits[40]),
    .S0N(ConfigBits_N[40]),
    .S1(ConfigBits[41]),
    .S1N(ConfigBits_N[41]),
    .X(J2MID_CDb_BEG0)
);
// switch matrix multiplexer J2MID_CDb_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDb_BEG1 (
    .A0(W2MID3),
    .A1(S2MID3),
    .A2(N2MID3),
    .A3(E2MID3),
    .S0(ConfigBits[42]),
    .S0N(ConfigBits_N[42]),
    .S1(ConfigBits[43]),
    .S1N(ConfigBits_N[43]),
    .X(J2MID_CDb_BEG1)
);
// switch matrix multiplexer J2MID_CDb_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDb_BEG2 (
    .A0(W2MID5),
    .A1(S2MID5),
    .A2(N2MID5),
    .A3(E2MID5),
    .S0(ConfigBits[44]),
    .S0N(ConfigBits_N[44]),
    .S1(ConfigBits[45]),
    .S1N(ConfigBits_N[45]),
    .X(J2MID_CDb_BEG2)
);
// switch matrix multiplexer J2MID_CDb_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_CDb_BEG3 (
    .A0(W2MID1),
    .A1(S2MID1),
    .A2(N2MID1),
    .A3(E2MID1),
    .S0(ConfigBits[46]),
    .S0N(ConfigBits_N[46]),
    .S1(ConfigBits[47]),
    .S1N(ConfigBits_N[47]),
    .X(J2MID_CDb_BEG3)
);
// switch matrix multiplexer J2MID_EFb_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFb_BEG0 (
    .A0(W2MID7),
    .A1(S2MID7),
    .A2(N2MID7),
    .A3(E2MID7),
    .S0(ConfigBits[48]),
    .S0N(ConfigBits_N[48]),
    .S1(ConfigBits[49]),
    .S1N(ConfigBits_N[49]),
    .X(J2MID_EFb_BEG0)
);
// switch matrix multiplexer J2MID_EFb_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFb_BEG1 (
    .A0(W2MID3),
    .A1(S2MID3),
    .A2(N2MID3),
    .A3(E2MID3),
    .S0(ConfigBits[50]),
    .S0N(ConfigBits_N[50]),
    .S1(ConfigBits[51]),
    .S1N(ConfigBits_N[51]),
    .X(J2MID_EFb_BEG1)
);
// switch matrix multiplexer J2MID_EFb_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFb_BEG2 (
    .A0(W2MID5),
    .A1(S2MID5),
    .A2(N2MID5),
    .A3(E2MID5),
    .S0(ConfigBits[52]),
    .S0N(ConfigBits_N[52]),
    .S1(ConfigBits[53]),
    .S1N(ConfigBits_N[53]),
    .X(J2MID_EFb_BEG2)
);
// switch matrix multiplexer J2MID_EFb_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_EFb_BEG3 (
    .A0(W2MID1),
    .A1(S2MID1),
    .A2(N2MID1),
    .A3(E2MID1),
    .S0(ConfigBits[54]),
    .S0N(ConfigBits_N[54]),
    .S1(ConfigBits[55]),
    .S1N(ConfigBits_N[55]),
    .X(J2MID_EFb_BEG3)
);
// switch matrix multiplexer J2MID_GHb_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHb_BEG0 (
    .A0(W2MID7),
    .A1(S2MID7),
    .A2(N2MID7),
    .A3(E2MID7),
    .S0(ConfigBits[56]),
    .S0N(ConfigBits_N[56]),
    .S1(ConfigBits[57]),
    .S1N(ConfigBits_N[57]),
    .X(J2MID_GHb_BEG0)
);
// switch matrix multiplexer J2MID_GHb_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHb_BEG1 (
    .A0(W2MID3),
    .A1(S2MID3),
    .A2(N2MID3),
    .A3(E2MID3),
    .S0(ConfigBits[58]),
    .S0N(ConfigBits_N[58]),
    .S1(ConfigBits[59]),
    .S1N(ConfigBits_N[59]),
    .X(J2MID_GHb_BEG1)
);
// switch matrix multiplexer J2MID_GHb_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHb_BEG2 (
    .A0(W2MID5),
    .A1(S2MID5),
    .A2(N2MID5),
    .A3(E2MID5),
    .S0(ConfigBits[60]),
    .S0N(ConfigBits_N[60]),
    .S1(ConfigBits[61]),
    .S1N(ConfigBits_N[61]),
    .X(J2MID_GHb_BEG2)
);
// switch matrix multiplexer J2MID_GHb_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2MID_GHb_BEG3 (
    .A0(W2MID1),
    .A1(S2MID1),
    .A2(N2MID1),
    .A3(E2MID1),
    .S0(ConfigBits[62]),
    .S0N(ConfigBits_N[62]),
    .S1(ConfigBits[63]),
    .S1N(ConfigBits_N[63]),
    .X(J2MID_GHb_BEG3)
);
// switch matrix multiplexer J2END_AB_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_AB_BEG0 (
    .A0(W2END6),
    .A1(SS4END3),
    .A2(N2END6),
    .A3(E2END6),
    .S0(ConfigBits[64]),
    .S0N(ConfigBits_N[64]),
    .S1(ConfigBits[65]),
    .S1N(ConfigBits_N[65]),
    .X(J2END_AB_BEG0)
);
// switch matrix multiplexer J2END_AB_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_AB_BEG1 (
    .A0(W2END2),
    .A1(S2END2),
    .A2(NN4END0),
    .A3(E2END2),
    .S0(ConfigBits[66]),
    .S0N(ConfigBits_N[66]),
    .S1(ConfigBits[67]),
    .S1N(ConfigBits_N[67]),
    .X(J2END_AB_BEG1)
);
// switch matrix multiplexer J2END_AB_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_AB_BEG2 (
    .A0(W2END4),
    .A1(S2END4),
    .A2(N2END4),
    .A3(EE4END0),
    .S0(ConfigBits[68]),
    .S0N(ConfigBits_N[68]),
    .S1(ConfigBits[69]),
    .S1N(ConfigBits_N[69]),
    .X(J2END_AB_BEG2)
);
// switch matrix multiplexer J2END_AB_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_AB_BEG3 (
    .A0(WW4END3),
    .A1(S2END0),
    .A2(N2END0),
    .A3(E2END0),
    .S0(ConfigBits[70]),
    .S0N(ConfigBits_N[70]),
    .S1(ConfigBits[71]),
    .S1N(ConfigBits_N[71]),
    .X(J2END_AB_BEG3)
);
// switch matrix multiplexer J2END_CD_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_CD_BEG0 (
    .A0(W2END6),
    .A1(S2END6),
    .A2(NN4END3),
    .A3(E2END6),
    .S0(ConfigBits[72]),
    .S0N(ConfigBits_N[72]),
    .S1(ConfigBits[73]),
    .S1N(ConfigBits_N[73]),
    .X(J2END_CD_BEG0)
);
// switch matrix multiplexer J2END_CD_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_CD_BEG1 (
    .A0(WW4END2),
    .A1(S2END2),
    .A2(N2END2),
    .A3(E2END2),
    .S0(ConfigBits[74]),
    .S0N(ConfigBits_N[74]),
    .S1(ConfigBits[75]),
    .S1N(ConfigBits_N[75]),
    .X(J2END_CD_BEG1)
);
// switch matrix multiplexer J2END_CD_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_CD_BEG2 (
    .A0(W2END4),
    .A1(SS4END2),
    .A2(N2END4),
    .A3(E2END4),
    .S0(ConfigBits[76]),
    .S0N(ConfigBits_N[76]),
    .S1(ConfigBits[77]),
    .S1N(ConfigBits_N[77]),
    .X(J2END_CD_BEG2)
);
// switch matrix multiplexer J2END_CD_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_CD_BEG3 (
    .A0(W2END0),
    .A1(S2END0),
    .A2(N2END0),
    .A3(EE4END1),
    .S0(ConfigBits[78]),
    .S0N(ConfigBits_N[78]),
    .S1(ConfigBits[79]),
    .S1N(ConfigBits_N[79]),
    .X(J2END_CD_BEG3)
);
// switch matrix multiplexer J2END_EF_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_EF_BEG0 (
    .A0(W2END7),
    .A1(S2END7),
    .A2(N2END7),
    .A3(EE4END2),
    .S0(ConfigBits[80]),
    .S0N(ConfigBits_N[80]),
    .S1(ConfigBits[81]),
    .S1N(ConfigBits_N[81]),
    .X(J2END_EF_BEG0)
);
// switch matrix multiplexer J2END_EF_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_EF_BEG1 (
    .A0(WW4END1),
    .A1(S2END3),
    .A2(N2END3),
    .A3(E2END3),
    .S0(ConfigBits[82]),
    .S0N(ConfigBits_N[82]),
    .S1(ConfigBits[83]),
    .S1N(ConfigBits_N[83]),
    .X(J2END_EF_BEG1)
);
// switch matrix multiplexer J2END_EF_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_EF_BEG2 (
    .A0(W2END5),
    .A1(SS4END1),
    .A2(N2END5),
    .A3(E2END5),
    .S0(ConfigBits[84]),
    .S0N(ConfigBits_N[84]),
    .S1(ConfigBits[85]),
    .S1N(ConfigBits_N[85]),
    .X(J2END_EF_BEG2)
);
// switch matrix multiplexer J2END_EF_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_EF_BEG3 (
    .A0(W2END1),
    .A1(S2END1),
    .A2(NN4END2),
    .A3(E2END1),
    .S0(ConfigBits[86]),
    .S0N(ConfigBits_N[86]),
    .S1(ConfigBits[87]),
    .S1N(ConfigBits_N[87]),
    .X(J2END_EF_BEG3)
);
// switch matrix multiplexer J2END_GH_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_GH_BEG0 (
    .A0(WW4END0),
    .A1(S2END7),
    .A2(N2END7),
    .A3(E2END7),
    .S0(ConfigBits[88]),
    .S0N(ConfigBits_N[88]),
    .S1(ConfigBits[89]),
    .S1N(ConfigBits_N[89]),
    .X(J2END_GH_BEG0)
);
// switch matrix multiplexer J2END_GH_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_GH_BEG1 (
    .A0(W2END3),
    .A1(SS4END0),
    .A2(N2END3),
    .A3(E2END3),
    .S0(ConfigBits[90]),
    .S0N(ConfigBits_N[90]),
    .S1(ConfigBits[91]),
    .S1N(ConfigBits_N[91]),
    .X(J2END_GH_BEG1)
);
// switch matrix multiplexer J2END_GH_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_GH_BEG2 (
    .A0(W2END5),
    .A1(S2END5),
    .A2(NN4END1),
    .A3(E2END5),
    .S0(ConfigBits[92]),
    .S0N(ConfigBits_N[92]),
    .S1(ConfigBits[93]),
    .S1N(ConfigBits_N[93]),
    .X(J2END_GH_BEG2)
);
// switch matrix multiplexer J2END_GH_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J2END_GH_BEG3 (
    .A0(W2END1),
    .A1(S2END1),
    .A2(N2END1),
    .A3(EE4END3),
    .S0(ConfigBits[94]),
    .S0N(ConfigBits_N[94]),
    .S1(ConfigBits[95]),
    .S1N(ConfigBits_N[95]),
    .X(J2END_GH_BEG3)
);
// switch matrix multiplexer J_l_AB_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_AB_BEG0 (
    .A0(WW4END0),
    .A1(S4END3),
    .A2(NN4END3),
    .A3(JN2END1),
    .S0(ConfigBits[96]),
    .S0N(ConfigBits_N[96]),
    .S1(ConfigBits[97]),
    .S1N(ConfigBits_N[97]),
    .X(J_l_AB_BEG0)
);
// switch matrix multiplexer J_l_AB_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_AB_BEG1 (
    .A0(W2END7),
    .A1(S4END2),
    .A2(JE2END1),
    .A3(EE4END2),
    .S0(ConfigBits[98]),
    .S0N(ConfigBits_N[98]),
    .S1(ConfigBits[99]),
    .S1N(ConfigBits_N[99]),
    .X(J_l_AB_BEG1)
);
// switch matrix multiplexer J_l_AB_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_AB_BEG2 (
    .A0(W6END1),
    .A1(JS2END1),
    .A2(N4END1),
    .A3(E6END1),
    .S0(ConfigBits[100]),
    .S0N(ConfigBits_N[100]),
    .S1(ConfigBits[101]),
    .S1N(ConfigBits_N[101]),
    .X(J_l_AB_BEG2)
);
// switch matrix multiplexer J_l_AB_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_AB_BEG3 (
    .A0(JW2END1),
    .A1(S4END0),
    .A2(N4END0),
    .A3(E6END0),
    .S0(ConfigBits[102]),
    .S0N(ConfigBits_N[102]),
    .S1(ConfigBits[103]),
    .S1N(ConfigBits_N[103]),
    .X(J_l_AB_BEG3)
);
// switch matrix multiplexer J_l_CD_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_CD_BEG0 (
    .A0(WW4END2),
    .A1(SS4END3),
    .A2(JN2END2),
    .A3(E2END3),
    .S0(ConfigBits[104]),
    .S0N(ConfigBits_N[104]),
    .S1(ConfigBits[105]),
    .S1N(ConfigBits_N[105]),
    .X(J_l_CD_BEG0)
);
// switch matrix multiplexer J_l_CD_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_CD_BEG1 (
    .A0(W2END7),
    .A1(JE2END2),
    .A2(N4END2),
    .A3(E2END2),
    .S0(ConfigBits[106]),
    .S0N(ConfigBits_N[106]),
    .S1(ConfigBits[107]),
    .S1N(ConfigBits_N[107]),
    .X(J_l_CD_BEG1)
);
// switch matrix multiplexer J_l_CD_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_CD_BEG2 (
    .A0(JS2END2),
    .A1(S4END1),
    .A2(NN4END1),
    .A3(EE4END1),
    .S0(ConfigBits[108]),
    .S0N(ConfigBits_N[108]),
    .S1(ConfigBits[109]),
    .S1N(ConfigBits_N[109]),
    .X(J_l_CD_BEG2)
);
// switch matrix multiplexer J_l_CD_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_CD_BEG3 (
    .A0(W6END0),
    .A1(SS4END0),
    .A2(N4END0),
    .A3(JW2END2),
    .S0(ConfigBits[110]),
    .S0N(ConfigBits_N[110]),
    .S1(ConfigBits[111]),
    .S1N(ConfigBits_N[111]),
    .X(J_l_CD_BEG3)
);
// switch matrix multiplexer J_l_EF_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_EF_BEG0 (
    .A0(W2END3),
    .A1(JN2END3),
    .A2(N4END3),
    .A3(E2END3),
    .S0(ConfigBits[112]),
    .S0N(ConfigBits_N[112]),
    .S1(ConfigBits[113]),
    .S1N(ConfigBits_N[113]),
    .X(J_l_EF_BEG0)
);
// switch matrix multiplexer J_l_EF_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_EF_BEG1 (
    .A0(JE2END3),
    .A1(S4END2),
    .A2(NN4END2),
    .A3(E2END2),
    .S0(ConfigBits[114]),
    .S0N(ConfigBits_N[114]),
    .S1(ConfigBits[115]),
    .S1N(ConfigBits_N[115]),
    .X(J_l_EF_BEG1)
);
// switch matrix multiplexer J_l_EF_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_EF_BEG2 (
    .A0(W2END4),
    .A1(SS4END1),
    .A2(N4END1),
    .A3(JS2END3),
    .S0(ConfigBits[116]),
    .S0N(ConfigBits_N[116]),
    .S1(ConfigBits[117]),
    .S1N(ConfigBits_N[117]),
    .X(J_l_EF_BEG2)
);
// switch matrix multiplexer J_l_EF_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_EF_BEG3 (
    .A0(WW4END1),
    .A1(S4END0),
    .A2(JW2END3),
    .A3(EE4END3),
    .S0(ConfigBits[118]),
    .S0N(ConfigBits_N[118]),
    .S1(ConfigBits[119]),
    .S1N(ConfigBits_N[119]),
    .X(J_l_EF_BEG3)
);
// switch matrix multiplexer J_l_GH_BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_GH_BEG0 (
    .A0(JN2END4),
    .A1(S4END3),
    .A2(N4END3),
    .A3(EE4END0),
    .S0(ConfigBits[120]),
    .S0N(ConfigBits_N[120]),
    .S1(ConfigBits[121]),
    .S1N(ConfigBits_N[121]),
    .X(J_l_GH_BEG0)
);
// switch matrix multiplexer J_l_GH_BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_GH_BEG1 (
    .A0(W2END2),
    .A1(SS4END2),
    .A2(N4END2),
    .A3(JE2END4),
    .S0(ConfigBits[122]),
    .S0N(ConfigBits_N[122]),
    .S1(ConfigBits[123]),
    .S1N(ConfigBits_N[123]),
    .X(J_l_GH_BEG1)
);
// switch matrix multiplexer J_l_GH_BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_GH_BEG2 (
    .A0(WW4END3),
    .A1(S4END1),
    .A2(JS2END4),
    .A3(E6END1),
    .S0(ConfigBits[124]),
    .S0N(ConfigBits_N[124]),
    .S1(ConfigBits[125]),
    .S1N(ConfigBits_N[125]),
    .X(J_l_GH_BEG2)
);
// switch matrix multiplexer J_l_GH_BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_J_l_GH_BEG3 (
    .A0(W2END0),
    .A1(JW2END4),
    .A2(NN4END0),
    .A3(E6END0),
    .S0(ConfigBits[126]),
    .S0N(ConfigBits_N[126]),
    .S1(ConfigBits[127]),
    .S1N(ConfigBits_N[127]),
    .X(J_l_GH_BEG3)
);
// switch matrix multiplexer LA_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LA_I0 (
    .A0(J_l_AB_END0),
    .A1(J2END_AB_END0),
    .A2(J2MID_ABb_END0),
    .A3(J2MID_ABa_END0),
    .S0(ConfigBits[128]),
    .S0N(ConfigBits_N[128]),
    .S1(ConfigBits[129]),
    .S1N(ConfigBits_N[129]),
    .X(LA_I0)
);
// switch matrix multiplexer LB_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LB_I0 (
    .A0(J_l_AB_END0),
    .A1(J2END_AB_END0),
    .A2(J2MID_ABb_END0),
    .A3(J2MID_ABa_END0),
    .S0(ConfigBits[130]),
    .S0N(ConfigBits_N[130]),
    .S1(ConfigBits[131]),
    .S1N(ConfigBits_N[131]),
    .X(LB_I0)
);
// switch matrix multiplexer LA_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LA_I1 (
    .A0(J_l_AB_END1),
    .A1(J2END_AB_END1),
    .A2(J2MID_ABb_END1),
    .A3(J2MID_ABa_END1),
    .S0(ConfigBits[132]),
    .S0N(ConfigBits_N[132]),
    .S1(ConfigBits[133]),
    .S1N(ConfigBits_N[133]),
    .X(LA_I1)
);
// switch matrix multiplexer LB_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LB_I1 (
    .A0(J_l_AB_END1),
    .A1(J2END_AB_END1),
    .A2(J2MID_ABb_END1),
    .A3(J2MID_ABa_END1),
    .S0(ConfigBits[134]),
    .S0N(ConfigBits_N[134]),
    .S1(ConfigBits[135]),
    .S1N(ConfigBits_N[135]),
    .X(LB_I1)
);
// switch matrix multiplexer LA_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LA_I2 (
    .A0(J_l_AB_END2),
    .A1(J2END_AB_END2),
    .A2(J2MID_ABb_END2),
    .A3(J2MID_ABa_END2),
    .S0(ConfigBits[136]),
    .S0N(ConfigBits_N[136]),
    .S1(ConfigBits[137]),
    .S1N(ConfigBits_N[137]),
    .X(LA_I2)
);
// switch matrix multiplexer LB_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LB_I2 (
    .A0(J_l_AB_END2),
    .A1(J2END_AB_END2),
    .A2(J2MID_ABb_END2),
    .A3(J2MID_ABa_END2),
    .S0(ConfigBits[138]),
    .S0N(ConfigBits_N[138]),
    .S1(ConfigBits[139]),
    .S1N(ConfigBits_N[139]),
    .X(LB_I2)
);
// switch matrix multiplexer LA_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LA_I3 (
    .A0(J_l_AB_END3),
    .A1(J2END_AB_END3),
    .A2(J2MID_ABb_END3),
    .A3(J2MID_ABa_END3),
    .S0(ConfigBits[140]),
    .S0N(ConfigBits_N[140]),
    .S1(ConfigBits[141]),
    .S1N(ConfigBits_N[141]),
    .X(LA_I3)
);
// switch matrix multiplexer LB_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LB_I3 (
    .A0(J_l_AB_END3),
    .A1(J2END_AB_END3),
    .A2(J2MID_ABb_END3),
    .A3(J2MID_ABa_END3),
    .S0(ConfigBits[142]),
    .S0N(ConfigBits_N[142]),
    .S1(ConfigBits[143]),
    .S1N(ConfigBits_N[143]),
    .X(LB_I3)
);
// switch matrix multiplexer LC_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LC_I0 (
    .A0(J_l_CD_END0),
    .A1(J2END_CD_END0),
    .A2(J2MID_CDb_END0),
    .A3(J2MID_CDa_END0),
    .S0(ConfigBits[144]),
    .S0N(ConfigBits_N[144]),
    .S1(ConfigBits[145]),
    .S1N(ConfigBits_N[145]),
    .X(LC_I0)
);
// switch matrix multiplexer LD_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LD_I0 (
    .A0(J_l_CD_END0),
    .A1(J2END_CD_END0),
    .A2(J2MID_CDb_END0),
    .A3(J2MID_CDa_END0),
    .S0(ConfigBits[146]),
    .S0N(ConfigBits_N[146]),
    .S1(ConfigBits[147]),
    .S1N(ConfigBits_N[147]),
    .X(LD_I0)
);
// switch matrix multiplexer LC_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LC_I1 (
    .A0(J_l_CD_END1),
    .A1(J2END_CD_END1),
    .A2(J2MID_CDb_END1),
    .A3(J2MID_CDa_END1),
    .S0(ConfigBits[148]),
    .S0N(ConfigBits_N[148]),
    .S1(ConfigBits[149]),
    .S1N(ConfigBits_N[149]),
    .X(LC_I1)
);
// switch matrix multiplexer LD_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LD_I1 (
    .A0(J_l_CD_END1),
    .A1(J2END_CD_END1),
    .A2(J2MID_CDb_END1),
    .A3(J2MID_CDa_END1),
    .S0(ConfigBits[150]),
    .S0N(ConfigBits_N[150]),
    .S1(ConfigBits[151]),
    .S1N(ConfigBits_N[151]),
    .X(LD_I1)
);
// switch matrix multiplexer LC_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LC_I2 (
    .A0(J_l_CD_END2),
    .A1(J2END_CD_END2),
    .A2(J2MID_CDb_END2),
    .A3(J2MID_CDa_END2),
    .S0(ConfigBits[152]),
    .S0N(ConfigBits_N[152]),
    .S1(ConfigBits[153]),
    .S1N(ConfigBits_N[153]),
    .X(LC_I2)
);
// switch matrix multiplexer LD_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LD_I2 (
    .A0(J_l_CD_END2),
    .A1(J2END_CD_END2),
    .A2(J2MID_CDb_END2),
    .A3(J2MID_CDa_END2),
    .S0(ConfigBits[154]),
    .S0N(ConfigBits_N[154]),
    .S1(ConfigBits[155]),
    .S1N(ConfigBits_N[155]),
    .X(LD_I2)
);
// switch matrix multiplexer LC_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LC_I3 (
    .A0(J_l_CD_END3),
    .A1(J2END_CD_END3),
    .A2(J2MID_CDb_END3),
    .A3(J2MID_CDa_END3),
    .S0(ConfigBits[156]),
    .S0N(ConfigBits_N[156]),
    .S1(ConfigBits[157]),
    .S1N(ConfigBits_N[157]),
    .X(LC_I3)
);
// switch matrix multiplexer LD_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LD_I3 (
    .A0(J_l_CD_END3),
    .A1(J2END_CD_END3),
    .A2(J2MID_CDb_END3),
    .A3(J2MID_CDa_END3),
    .S0(ConfigBits[158]),
    .S0N(ConfigBits_N[158]),
    .S1(ConfigBits[159]),
    .S1N(ConfigBits_N[159]),
    .X(LD_I3)
);
// switch matrix multiplexer LE_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LE_I0 (
    .A0(J_l_EF_END0),
    .A1(J2END_EF_END0),
    .A2(J2MID_EFb_END0),
    .A3(J2MID_EFa_END0),
    .S0(ConfigBits[160]),
    .S0N(ConfigBits_N[160]),
    .S1(ConfigBits[161]),
    .S1N(ConfigBits_N[161]),
    .X(LE_I0)
);
// switch matrix multiplexer LF_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LF_I0 (
    .A0(J_l_EF_END0),
    .A1(J2END_EF_END0),
    .A2(J2MID_EFb_END0),
    .A3(J2MID_EFa_END0),
    .S0(ConfigBits[162]),
    .S0N(ConfigBits_N[162]),
    .S1(ConfigBits[163]),
    .S1N(ConfigBits_N[163]),
    .X(LF_I0)
);
// switch matrix multiplexer LE_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LE_I1 (
    .A0(J_l_EF_END1),
    .A1(J2END_EF_END1),
    .A2(J2MID_EFb_END1),
    .A3(J2MID_EFa_END1),
    .S0(ConfigBits[164]),
    .S0N(ConfigBits_N[164]),
    .S1(ConfigBits[165]),
    .S1N(ConfigBits_N[165]),
    .X(LE_I1)
);
// switch matrix multiplexer LF_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LF_I1 (
    .A0(J_l_EF_END1),
    .A1(J2END_EF_END1),
    .A2(J2MID_EFb_END1),
    .A3(J2MID_EFa_END1),
    .S0(ConfigBits[166]),
    .S0N(ConfigBits_N[166]),
    .S1(ConfigBits[167]),
    .S1N(ConfigBits_N[167]),
    .X(LF_I1)
);
// switch matrix multiplexer LE_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LE_I2 (
    .A0(J_l_EF_END2),
    .A1(J2END_EF_END2),
    .A2(J2MID_EFb_END2),
    .A3(J2MID_EFa_END2),
    .S0(ConfigBits[168]),
    .S0N(ConfigBits_N[168]),
    .S1(ConfigBits[169]),
    .S1N(ConfigBits_N[169]),
    .X(LE_I2)
);
// switch matrix multiplexer LF_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LF_I2 (
    .A0(J_l_EF_END2),
    .A1(J2END_EF_END2),
    .A2(J2MID_EFb_END2),
    .A3(J2MID_EFa_END2),
    .S0(ConfigBits[170]),
    .S0N(ConfigBits_N[170]),
    .S1(ConfigBits[171]),
    .S1N(ConfigBits_N[171]),
    .X(LF_I2)
);
// switch matrix multiplexer LE_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LE_I3 (
    .A0(J_l_EF_END3),
    .A1(J2END_EF_END3),
    .A2(J2MID_EFb_END3),
    .A3(J2MID_EFa_END3),
    .S0(ConfigBits[172]),
    .S0N(ConfigBits_N[172]),
    .S1(ConfigBits[173]),
    .S1N(ConfigBits_N[173]),
    .X(LE_I3)
);
// switch matrix multiplexer LF_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LF_I3 (
    .A0(J_l_EF_END3),
    .A1(J2END_EF_END3),
    .A2(J2MID_EFb_END3),
    .A3(J2MID_EFa_END3),
    .S0(ConfigBits[174]),
    .S0N(ConfigBits_N[174]),
    .S1(ConfigBits[175]),
    .S1N(ConfigBits_N[175]),
    .X(LF_I3)
);
// switch matrix multiplexer LG_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LG_I0 (
    .A0(J_l_GH_END0),
    .A1(J2END_GH_END0),
    .A2(J2MID_GHb_END0),
    .A3(J2MID_GHa_END0),
    .S0(ConfigBits[176]),
    .S0N(ConfigBits_N[176]),
    .S1(ConfigBits[177]),
    .S1N(ConfigBits_N[177]),
    .X(LG_I0)
);
// switch matrix multiplexer LH_I0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LH_I0 (
    .A0(J_l_GH_END0),
    .A1(J2END_GH_END0),
    .A2(J2MID_GHb_END0),
    .A3(J2MID_GHa_END0),
    .S0(ConfigBits[178]),
    .S0N(ConfigBits_N[178]),
    .S1(ConfigBits[179]),
    .S1N(ConfigBits_N[179]),
    .X(LH_I0)
);
// switch matrix multiplexer LG_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LG_I1 (
    .A0(J_l_GH_END1),
    .A1(J2END_GH_END1),
    .A2(J2MID_GHb_END1),
    .A3(J2MID_GHa_END1),
    .S0(ConfigBits[180]),
    .S0N(ConfigBits_N[180]),
    .S1(ConfigBits[181]),
    .S1N(ConfigBits_N[181]),
    .X(LG_I1)
);
// switch matrix multiplexer LH_I1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LH_I1 (
    .A0(J_l_GH_END1),
    .A1(J2END_GH_END1),
    .A2(J2MID_GHb_END1),
    .A3(J2MID_GHa_END1),
    .S0(ConfigBits[182]),
    .S0N(ConfigBits_N[182]),
    .S1(ConfigBits[183]),
    .S1N(ConfigBits_N[183]),
    .X(LH_I1)
);
// switch matrix multiplexer LG_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LG_I2 (
    .A0(J_l_GH_END2),
    .A1(J2END_GH_END2),
    .A2(J2MID_GHb_END2),
    .A3(J2MID_GHa_END2),
    .S0(ConfigBits[184]),
    .S0N(ConfigBits_N[184]),
    .S1(ConfigBits[185]),
    .S1N(ConfigBits_N[185]),
    .X(LG_I2)
);
// switch matrix multiplexer LH_I2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LH_I2 (
    .A0(J_l_GH_END2),
    .A1(J2END_GH_END2),
    .A2(J2MID_GHb_END2),
    .A3(J2MID_GHa_END2),
    .S0(ConfigBits[186]),
    .S0N(ConfigBits_N[186]),
    .S1(ConfigBits[187]),
    .S1N(ConfigBits_N[187]),
    .X(LH_I2)
);
// switch matrix multiplexer LG_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LG_I3 (
    .A0(J_l_GH_END3),
    .A1(J2END_GH_END3),
    .A2(J2MID_GHb_END3),
    .A3(J2MID_GHa_END3),
    .S0(ConfigBits[188]),
    .S0N(ConfigBits_N[188]),
    .S1(ConfigBits[189]),
    .S1N(ConfigBits_N[189]),
    .X(LG_I3)
);
// switch matrix multiplexer LH_I3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_LH_I3 (
    .A0(J_l_GH_END3),
    .A1(J2END_GH_END3),
    .A2(J2MID_GHb_END3),
    .A3(J2MID_GHa_END3),
    .S0(ConfigBits[190]),
    .S0N(ConfigBits_N[190]),
    .S1(ConfigBits[191]),
    .S1N(ConfigBits_N[191]),
    .X(LH_I3)
);
// switch matrix multiplexer JN2BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG0 (
    .A0(N4END1),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END1),
    .A4(SS4END1),
    .A5(E2END1),
    .A6(N2END1),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(E1END3),
    .S0(ConfigBits[192]),
    .S0N(ConfigBits_N[192]),
    .S1(ConfigBits[193]),
    .S1N(ConfigBits_N[193]),
    .S2(ConfigBits[194]),
    .S2N(ConfigBits_N[194]),
    .S3(ConfigBits[195]),
    .S3N(ConfigBits_N[195]),
    .X(JN2BEG0)
);
// switch matrix multiplexer JN2BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG1 (
    .A0(N4END2),
    .A1(E6END0),
    .A2(W6END0),
    .A3(W2END2),
    .A4(S2END2),
    .A5(E2END2),
    .A6(N2END2),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(E1END0),
    .A15(LA_O),
    .S0(ConfigBits[196]),
    .S0N(ConfigBits_N[196]),
    .S1(ConfigBits[197]),
    .S1N(ConfigBits_N[197]),
    .S2(ConfigBits[198]),
    .S2N(ConfigBits_N[198]),
    .S3(ConfigBits[199]),
    .S3N(ConfigBits_N[199]),
    .X(JN2BEG1)
);
// switch matrix multiplexer JN2BEG2 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG2 (
    .A0(N4END3),
    .A1(E6END1),
    .A2(WW4END1),
    .A3(W2END3),
    .A4(S2END3),
    .A5(E2END3),
    .A6(N2END3),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(E1END1),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[200]),
    .S0N(ConfigBits_N[200]),
    .S1(ConfigBits[201]),
    .S1N(ConfigBits_N[201]),
    .S2(ConfigBits[202]),
    .S2N(ConfigBits_N[202]),
    .S3(ConfigBits[203]),
    .S3N(ConfigBits_N[203]),
    .X(JN2BEG2)
);
// switch matrix multiplexer JN2BEG3 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG3 (
    .A0(N4END0),
    .A1(E6END0),
    .A2(W6END0),
    .A3(W2END4),
    .A4(S2END4),
    .A5(E2END4),
    .A6(N2END4),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(E1END2),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[204]),
    .S0N(ConfigBits_N[204]),
    .S1(ConfigBits[205]),
    .S1N(ConfigBits_N[205]),
    .S2(ConfigBits[206]),
    .S2N(ConfigBits_N[206]),
    .S3(ConfigBits[207]),
    .S3N(ConfigBits_N[207]),
    .X(JN2BEG3)
);
// switch matrix multiplexer JN2BEG4 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG4 (
    .A0(W1END1),
    .A1(S1END1),
    .A2(E1END1),
    .A3(N1END1),
    .A4(S2END5),
    .A5(E2END5),
    .A6(N2END5),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(W1END3),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[208]),
    .S0N(ConfigBits_N[208]),
    .S1(ConfigBits[209]),
    .S1N(ConfigBits_N[209]),
    .S2(ConfigBits[210]),
    .S2N(ConfigBits_N[210]),
    .S3(ConfigBits[211]),
    .S3N(ConfigBits_N[211]),
    .X(JN2BEG4)
);
// switch matrix multiplexer JN2BEG5 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG5 (
    .A0(W1END2),
    .A1(S1END2),
    .A2(E1END2),
    .A3(N1END2),
    .A4(S2END6),
    .A5(E2END6),
    .A6(N2END6),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(W1END0),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[212]),
    .S0N(ConfigBits_N[212]),
    .S1(ConfigBits[213]),
    .S1N(ConfigBits_N[213]),
    .S2(ConfigBits[214]),
    .S2N(ConfigBits_N[214]),
    .S3(ConfigBits[215]),
    .S3N(ConfigBits_N[215]),
    .X(JN2BEG5)
);
// switch matrix multiplexer JN2BEG6 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG6 (
    .A0(W1END3),
    .A1(S1END3),
    .A2(E1END3),
    .A3(N1END3),
    .A4(S2END7),
    .A5(E2END7),
    .A6(N2END7),
    .A7(M_AH),
    .A8(LH_O),
    .A9(W1END1),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[216]),
    .S0N(ConfigBits_N[216]),
    .S1(ConfigBits[217]),
    .S1N(ConfigBits_N[217]),
    .S2(ConfigBits[218]),
    .S2N(ConfigBits_N[218]),
    .S3(ConfigBits[219]),
    .S3N(ConfigBits_N[219]),
    .X(JN2BEG6)
);
// switch matrix multiplexer JN2BEG7 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JN2BEG7 (
    .A0(W1END0),
    .A1(S1END0),
    .A2(E1END0),
    .A3(N1END0),
    .A4(S2END0),
    .A5(EE4END0),
    .A6(N2END0),
    .A7(M_EF),
    .A8(W1END2),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[220]),
    .S0N(ConfigBits_N[220]),
    .S1(ConfigBits[221]),
    .S1N(ConfigBits_N[221]),
    .S2(ConfigBits[222]),
    .S2N(ConfigBits_N[222]),
    .S3(ConfigBits[223]),
    .S3N(ConfigBits_N[223]),
    .X(JN2BEG7)
);
// switch matrix multiplexer JE2BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG0 (
    .A0(N4END1),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END1),
    .A4(S2END1),
    .A5(EE4END1),
    .A6(N2END1),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(N1END3),
    .S0(ConfigBits[224]),
    .S0N(ConfigBits_N[224]),
    .S1(ConfigBits[225]),
    .S1N(ConfigBits_N[225]),
    .S2(ConfigBits[226]),
    .S2N(ConfigBits_N[226]),
    .S3(ConfigBits[227]),
    .S3N(ConfigBits_N[227]),
    .X(JE2BEG0)
);
// switch matrix multiplexer JE2BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG1 (
    .A0(N4END2),
    .A1(E6END0),
    .A2(WW4END3),
    .A3(W2END2),
    .A4(S2END2),
    .A5(E2END2),
    .A6(N2END2),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(N1END0),
    .A15(LA_O),
    .S0(ConfigBits[228]),
    .S0N(ConfigBits_N[228]),
    .S1(ConfigBits[229]),
    .S1N(ConfigBits_N[229]),
    .S2(ConfigBits[230]),
    .S2N(ConfigBits_N[230]),
    .S3(ConfigBits[231]),
    .S3N(ConfigBits_N[231]),
    .X(JE2BEG1)
);
// switch matrix multiplexer JE2BEG2 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG2 (
    .A0(N4END3),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END3),
    .A4(S2END3),
    .A5(E2END3),
    .A6(N2END3),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(N1END1),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[232]),
    .S0N(ConfigBits_N[232]),
    .S1(ConfigBits[233]),
    .S1N(ConfigBits_N[233]),
    .S2(ConfigBits[234]),
    .S2N(ConfigBits_N[234]),
    .S3(ConfigBits[235]),
    .S3N(ConfigBits_N[235]),
    .X(JE2BEG2)
);
// switch matrix multiplexer JE2BEG3 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG3 (
    .A0(N4END0),
    .A1(E6END0),
    .A2(W6END0),
    .A3(W2END4),
    .A4(S2END4),
    .A5(E2END4),
    .A6(N2END4),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(N1END2),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[236]),
    .S0N(ConfigBits_N[236]),
    .S1(ConfigBits[237]),
    .S1N(ConfigBits_N[237]),
    .S2(ConfigBits[238]),
    .S2N(ConfigBits_N[238]),
    .S3(ConfigBits[239]),
    .S3N(ConfigBits_N[239]),
    .X(JE2BEG3)
);
// switch matrix multiplexer JE2BEG4 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG4 (
    .A0(W1END1),
    .A1(S1END1),
    .A2(E1END1),
    .A3(N1END1),
    .A4(S2END5),
    .A5(E2END5),
    .A6(N2END5),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(S1END3),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[240]),
    .S0N(ConfigBits_N[240]),
    .S1(ConfigBits[241]),
    .S1N(ConfigBits_N[241]),
    .S2(ConfigBits[242]),
    .S2N(ConfigBits_N[242]),
    .S3(ConfigBits[243]),
    .S3N(ConfigBits_N[243]),
    .X(JE2BEG4)
);
// switch matrix multiplexer JE2BEG5 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG5 (
    .A0(W1END2),
    .A1(S1END2),
    .A2(E1END2),
    .A3(N1END2),
    .A4(S2END6),
    .A5(E2END6),
    .A6(N2END6),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(S1END0),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[244]),
    .S0N(ConfigBits_N[244]),
    .S1(ConfigBits[245]),
    .S1N(ConfigBits_N[245]),
    .S2(ConfigBits[246]),
    .S2N(ConfigBits_N[246]),
    .S3(ConfigBits[247]),
    .S3N(ConfigBits_N[247]),
    .X(JE2BEG5)
);
// switch matrix multiplexer JE2BEG6 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG6 (
    .A0(W1END3),
    .A1(S1END3),
    .A2(E1END3),
    .A3(N1END3),
    .A4(S2END7),
    .A5(E2END7),
    .A6(N2END7),
    .A7(M_AD),
    .A8(LH_O),
    .A9(S1END1),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[248]),
    .S0N(ConfigBits_N[248]),
    .S1(ConfigBits[249]),
    .S1N(ConfigBits_N[249]),
    .S2(ConfigBits[250]),
    .S2N(ConfigBits_N[250]),
    .S3(ConfigBits[251]),
    .S3N(ConfigBits_N[251]),
    .X(JE2BEG6)
);
// switch matrix multiplexer JE2BEG7 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JE2BEG7 (
    .A0(WW4END0),
    .A1(S1END0),
    .A2(E1END0),
    .A3(N1END0),
    .A4(SS4END0),
    .A5(E2END0),
    .A6(N2END0),
    .A7(M_AH),
    .A8(S1END2),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[252]),
    .S0N(ConfigBits_N[252]),
    .S1(ConfigBits[253]),
    .S1N(ConfigBits_N[253]),
    .S2(ConfigBits[254]),
    .S2N(ConfigBits_N[254]),
    .S3(ConfigBits[255]),
    .S3N(ConfigBits_N[255]),
    .X(JE2BEG7)
);
// switch matrix multiplexer JS2BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG0 (
    .A0(S4END1),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END1),
    .A4(S2END1),
    .A5(E2END1),
    .A6(NN4END1),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(E1END3),
    .S0(ConfigBits[256]),
    .S0N(ConfigBits_N[256]),
    .S1(ConfigBits[257]),
    .S1N(ConfigBits_N[257]),
    .S2(ConfigBits[258]),
    .S2N(ConfigBits_N[258]),
    .S3(ConfigBits[259]),
    .S3N(ConfigBits_N[259]),
    .X(JS2BEG0)
);
// switch matrix multiplexer JS2BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG1 (
    .A0(S4END2),
    .A1(E6END0),
    .A2(W6END0),
    .A3(W2END2),
    .A4(SS4END2),
    .A5(EE4END2),
    .A6(NN4END2),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(E1END0),
    .A15(LA_O),
    .S0(ConfigBits[260]),
    .S0N(ConfigBits_N[260]),
    .S1(ConfigBits[261]),
    .S1N(ConfigBits_N[261]),
    .S2(ConfigBits[262]),
    .S2N(ConfigBits_N[262]),
    .S3(ConfigBits[263]),
    .S3N(ConfigBits_N[263]),
    .X(JS2BEG1)
);
// switch matrix multiplexer JS2BEG2 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG2 (
    .A0(S4END3),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END3),
    .A4(S2END3),
    .A5(E2END3),
    .A6(NN4END3),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(E1END1),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[264]),
    .S0N(ConfigBits_N[264]),
    .S1(ConfigBits[265]),
    .S1N(ConfigBits_N[265]),
    .S2(ConfigBits[266]),
    .S2N(ConfigBits_N[266]),
    .S3(ConfigBits[267]),
    .S3N(ConfigBits_N[267]),
    .X(JS2BEG2)
);
// switch matrix multiplexer JS2BEG3 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG3 (
    .A0(S4END0),
    .A1(E6END0),
    .A2(WW4END2),
    .A3(W2END4),
    .A4(S2END4),
    .A5(E2END4),
    .A6(N2END4),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(E1END2),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[268]),
    .S0N(ConfigBits_N[268]),
    .S1(ConfigBits[269]),
    .S1N(ConfigBits_N[269]),
    .S2(ConfigBits[270]),
    .S2N(ConfigBits_N[270]),
    .S3(ConfigBits[271]),
    .S3N(ConfigBits_N[271]),
    .X(JS2BEG3)
);
// switch matrix multiplexer JS2BEG4 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG4 (
    .A0(W1END1),
    .A1(S1END1),
    .A2(E1END1),
    .A3(N1END1),
    .A4(S2END5),
    .A5(E2END5),
    .A6(N2END5),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(W1END3),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[272]),
    .S0N(ConfigBits_N[272]),
    .S1(ConfigBits[273]),
    .S1N(ConfigBits_N[273]),
    .S2(ConfigBits[274]),
    .S2N(ConfigBits_N[274]),
    .S3(ConfigBits[275]),
    .S3N(ConfigBits_N[275]),
    .X(JS2BEG4)
);
// switch matrix multiplexer JS2BEG5 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG5 (
    .A0(W1END2),
    .A1(S1END2),
    .A2(E1END2),
    .A3(N1END2),
    .A4(S2END6),
    .A5(E2END6),
    .A6(N2END6),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(W1END0),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[276]),
    .S0N(ConfigBits_N[276]),
    .S1(ConfigBits[277]),
    .S1N(ConfigBits_N[277]),
    .S2(ConfigBits[278]),
    .S2N(ConfigBits_N[278]),
    .S3(ConfigBits[279]),
    .S3N(ConfigBits_N[279]),
    .X(JS2BEG5)
);
// switch matrix multiplexer JS2BEG6 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG6 (
    .A0(W1END3),
    .A1(S1END3),
    .A2(E1END3),
    .A3(N1END3),
    .A4(S2END7),
    .A5(E2END7),
    .A6(N2END7),
    .A7(M_AB),
    .A8(LH_O),
    .A9(W1END1),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[280]),
    .S0N(ConfigBits_N[280]),
    .S1(ConfigBits[281]),
    .S1N(ConfigBits_N[281]),
    .S2(ConfigBits[282]),
    .S2N(ConfigBits_N[282]),
    .S3(ConfigBits[283]),
    .S3N(ConfigBits_N[283]),
    .X(JS2BEG6)
);
// switch matrix multiplexer JS2BEG7 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JS2BEG7 (
    .A0(W1END0),
    .A1(S1END0),
    .A2(E1END0),
    .A3(N1END0),
    .A4(S2END0),
    .A5(E2END0),
    .A6(N2END0),
    .A7(M_AD),
    .A8(W1END2),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[284]),
    .S0N(ConfigBits_N[284]),
    .S1(ConfigBits[285]),
    .S1N(ConfigBits_N[285]),
    .S2(ConfigBits[286]),
    .S2N(ConfigBits_N[286]),
    .S3(ConfigBits[287]),
    .S3N(ConfigBits_N[287]),
    .X(JS2BEG7)
);
// switch matrix multiplexer JW2BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG0 (
    .A0(S4END1),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END1),
    .A4(S2END1),
    .A5(E2END1),
    .A6(N2END1),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(N1END3),
    .S0(ConfigBits[288]),
    .S0N(ConfigBits_N[288]),
    .S1(ConfigBits[289]),
    .S1N(ConfigBits_N[289]),
    .S2(ConfigBits[290]),
    .S2N(ConfigBits_N[290]),
    .S3(ConfigBits[291]),
    .S3N(ConfigBits_N[291]),
    .X(JW2BEG0)
);
// switch matrix multiplexer JW2BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG1 (
    .A0(S4END2),
    .A1(E6END0),
    .A2(W6END0),
    .A3(W2END2),
    .A4(S2END2),
    .A5(E2END2),
    .A6(N2END2),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(N1END0),
    .A15(LA_O),
    .S0(ConfigBits[292]),
    .S0N(ConfigBits_N[292]),
    .S1(ConfigBits[293]),
    .S1N(ConfigBits_N[293]),
    .S2(ConfigBits[294]),
    .S2N(ConfigBits_N[294]),
    .S3(ConfigBits[295]),
    .S3N(ConfigBits_N[295]),
    .X(JW2BEG1)
);
// switch matrix multiplexer JW2BEG2 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG2 (
    .A0(S4END3),
    .A1(E6END1),
    .A2(W6END1),
    .A3(W2END3),
    .A4(SS4END3),
    .A5(EE4END3),
    .A6(N2END3),
    .A7(M_EF),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(N1END1),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[296]),
    .S0N(ConfigBits_N[296]),
    .S1(ConfigBits[297]),
    .S1N(ConfigBits_N[297]),
    .S2(ConfigBits[298]),
    .S2N(ConfigBits_N[298]),
    .S3(ConfigBits[299]),
    .S3N(ConfigBits_N[299]),
    .X(JW2BEG2)
);
// switch matrix multiplexer JW2BEG3 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG3 (
    .A0(S4END0),
    .A1(E6END0),
    .A2(WW4END2),
    .A3(W2END4),
    .A4(S2END4),
    .A5(E2END4),
    .A6(N2END4),
    .A7(M_AB),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(N1END2),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[300]),
    .S0N(ConfigBits_N[300]),
    .S1(ConfigBits[301]),
    .S1N(ConfigBits_N[301]),
    .S2(ConfigBits[302]),
    .S2N(ConfigBits_N[302]),
    .S3(ConfigBits[303]),
    .S3N(ConfigBits_N[303]),
    .X(JW2BEG3)
);
// switch matrix multiplexer JW2BEG4 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG4 (
    .A0(W1END1),
    .A1(S1END1),
    .A2(E1END1),
    .A3(N1END1),
    .A4(S2END5),
    .A5(E2END5),
    .A6(N2END5),
    .A7(M_AD),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(S1END3),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[304]),
    .S0N(ConfigBits_N[304]),
    .S1(ConfigBits[305]),
    .S1N(ConfigBits_N[305]),
    .S2(ConfigBits[306]),
    .S2N(ConfigBits_N[306]),
    .S3(ConfigBits[307]),
    .S3N(ConfigBits_N[307]),
    .X(JW2BEG4)
);
// switch matrix multiplexer JW2BEG5 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG5 (
    .A0(W1END2),
    .A1(S1END2),
    .A2(E1END2),
    .A3(N1END2),
    .A4(S2END6),
    .A5(E2END6),
    .A6(N2END6),
    .A7(M_AH),
    .A8(LH_O),
    .A9(LG_O),
    .A10(S1END0),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[308]),
    .S0N(ConfigBits_N[308]),
    .S1(ConfigBits[309]),
    .S1N(ConfigBits_N[309]),
    .S2(ConfigBits[310]),
    .S2N(ConfigBits_N[310]),
    .S3(ConfigBits[311]),
    .S3N(ConfigBits_N[311]),
    .X(JW2BEG5)
);
// switch matrix multiplexer JW2BEG6 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG6 (
    .A0(W1END3),
    .A1(S1END3),
    .A2(E1END3),
    .A3(N1END3),
    .A4(S2END7),
    .A5(E2END7),
    .A6(N2END7),
    .A7(M_EF),
    .A8(LH_O),
    .A9(S1END1),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[312]),
    .S0N(ConfigBits_N[312]),
    .S1(ConfigBits[313]),
    .S1N(ConfigBits_N[313]),
    .S2(ConfigBits[314]),
    .S2N(ConfigBits_N[314]),
    .S3(ConfigBits[315]),
    .S3N(ConfigBits_N[315]),
    .X(JW2BEG6)
);
// switch matrix multiplexer JW2BEG7 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_JW2BEG7 (
    .A0(W1END0),
    .A1(S1END0),
    .A2(E1END0),
    .A3(N1END0),
    .A4(S2END0),
    .A5(E2END0),
    .A6(NN4END0),
    .A7(M_AB),
    .A8(S1END2),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[316]),
    .S0N(ConfigBits_N[316]),
    .S1(ConfigBits[317]),
    .S1N(ConfigBits_N[317]),
    .S2(ConfigBits[318]),
    .S2N(ConfigBits_N[318]),
    .S3(ConfigBits[319]),
    .S3N(ConfigBits_N[319]),
    .X(JW2BEG7)
);
// switch matrix multiplexer N2BEG0 MUX-1assign N2BEG0 = JN2END0;// switch matrix multiplexer N2BEG1 MUX-1assign N2BEG1 = JN2END1;// switch matrix multiplexer N2BEG2 MUX-1assign N2BEG2 = JN2END2;// switch matrix multiplexer N2BEG3 MUX-1assign N2BEG3 = JN2END3;// switch matrix multiplexer N2BEG4 MUX-1assign N2BEG4 = JN2END4;// switch matrix multiplexer N2BEG5 MUX-1assign N2BEG5 = JN2END5;// switch matrix multiplexer N2BEG6 MUX-1assign N2BEG6 = JN2END6;// switch matrix multiplexer N2BEG7 MUX-1assign N2BEG7 = JN2END7;// switch matrix multiplexer E2BEG0 MUX-1assign E2BEG0 = JE2END0;// switch matrix multiplexer E2BEG1 MUX-1assign E2BEG1 = JE2END1;// switch matrix multiplexer E2BEG2 MUX-1assign E2BEG2 = JE2END2;// switch matrix multiplexer E2BEG3 MUX-1assign E2BEG3 = JE2END3;// switch matrix multiplexer E2BEG4 MUX-1assign E2BEG4 = JE2END4;// switch matrix multiplexer E2BEG5 MUX-1assign E2BEG5 = JE2END5;// switch matrix multiplexer E2BEG6 MUX-1assign E2BEG6 = JE2END6;// switch matrix multiplexer E2BEG7 MUX-1assign E2BEG7 = JE2END7;// switch matrix multiplexer S2BEG0 MUX-1assign S2BEG0 = JS2END0;// switch matrix multiplexer S2BEG1 MUX-1assign S2BEG1 = JS2END1;// switch matrix multiplexer S2BEG2 MUX-1assign S2BEG2 = JS2END2;// switch matrix multiplexer S2BEG3 MUX-1assign S2BEG3 = JS2END3;// switch matrix multiplexer S2BEG4 MUX-1assign S2BEG4 = JS2END4;// switch matrix multiplexer S2BEG5 MUX-1assign S2BEG5 = JS2END5;// switch matrix multiplexer S2BEG6 MUX-1assign S2BEG6 = JS2END6;// switch matrix multiplexer S2BEG7 MUX-1assign S2BEG7 = JS2END7;// switch matrix multiplexer W2BEG1 MUX-1assign W2BEG1 = JW2END1;// switch matrix multiplexer W2BEG2 MUX-1assign W2BEG2 = JW2END2;// switch matrix multiplexer W2BEG5 MUX-1assign W2BEG5 = JW2END5;// switch matrix multiplexer W2BEG6 MUX-1assign W2BEG6 = JW2END6;// switch matrix multiplexer W2BEG0 MUX-1assign W2BEG0 = JW2END0;// switch matrix multiplexer W2BEG3 MUX-1assign W2BEG3 = JW2END3;// switch matrix multiplexer W2BEG4 MUX-1assign W2BEG4 = JW2END4;// switch matrix multiplexer W2BEG7 MUX-1assign W2BEG7 = JW2END7;// switch matrix multiplexer N1BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N1BEG0 (
    .A0(J2MID_CDb_END3),
    .A1(JW2END3),
    .A2(LC_O),
    .A3(J_l_CD_END1),
    .S0(ConfigBits[320]),
    .S0N(ConfigBits_N[320]),
    .S1(ConfigBits[321]),
    .S1N(ConfigBits_N[321]),
    .X(N1BEG0)
);
// switch matrix multiplexer N1BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N1BEG1 (
    .A0(J2MID_EFb_END0),
    .A1(JW2END0),
    .A2(LD_O),
    .A3(J_l_EF_END2),
    .S0(ConfigBits[322]),
    .S0N(ConfigBits_N[322]),
    .S1(ConfigBits[323]),
    .S1N(ConfigBits_N[323]),
    .X(N1BEG1)
);
// switch matrix multiplexer N1BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N1BEG2 (
    .A0(J2MID_GHb_END1),
    .A1(JW2END1),
    .A2(LE_O),
    .A3(J_l_GH_END3),
    .S0(ConfigBits[324]),
    .S0N(ConfigBits_N[324]),
    .S1(ConfigBits[325]),
    .S1N(ConfigBits_N[325]),
    .X(N1BEG2)
);
// switch matrix multiplexer N1BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N1BEG3 (
    .A0(J2MID_ABb_END2),
    .A1(JW2END2),
    .A2(LF_O),
    .A3(J_l_AB_END0),
    .S0(ConfigBits[326]),
    .S0N(ConfigBits_N[326]),
    .S1(ConfigBits[327]),
    .S1N(ConfigBits_N[327]),
    .X(N1BEG3)
);
// switch matrix multiplexer E1BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_E1BEG0 (
    .A0(J2MID_CDb_END3),
    .A1(JN2END3),
    .A2(LD_O),
    .A3(J_l_CD_END1),
    .S0(ConfigBits[328]),
    .S0N(ConfigBits_N[328]),
    .S1(ConfigBits[329]),
    .S1N(ConfigBits_N[329]),
    .X(E1BEG0)
);
// switch matrix multiplexer E1BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_E1BEG1 (
    .A0(J2MID_EFb_END0),
    .A1(JN2END0),
    .A2(LE_O),
    .A3(J_l_EF_END2),
    .S0(ConfigBits[330]),
    .S0N(ConfigBits_N[330]),
    .S1(ConfigBits[331]),
    .S1N(ConfigBits_N[331]),
    .X(E1BEG1)
);
// switch matrix multiplexer E1BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_E1BEG2 (
    .A0(J2MID_GHb_END1),
    .A1(JN2END1),
    .A2(LF_O),
    .A3(J_l_GH_END3),
    .S0(ConfigBits[332]),
    .S0N(ConfigBits_N[332]),
    .S1(ConfigBits[333]),
    .S1N(ConfigBits_N[333]),
    .X(E1BEG2)
);
// switch matrix multiplexer E1BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_E1BEG3 (
    .A0(J2MID_ABb_END2),
    .A1(JN2END2),
    .A2(LG_O),
    .A3(J_l_AB_END0),
    .S0(ConfigBits[334]),
    .S0N(ConfigBits_N[334]),
    .S1(ConfigBits[335]),
    .S1N(ConfigBits_N[335]),
    .X(E1BEG3)
);
// switch matrix multiplexer S1BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S1BEG0 (
    .A0(J2MID_CDb_END3),
    .A1(JE2END3),
    .A2(LE_O),
    .A3(J_l_CD_END1),
    .S0(ConfigBits[336]),
    .S0N(ConfigBits_N[336]),
    .S1(ConfigBits[337]),
    .S1N(ConfigBits_N[337]),
    .X(S1BEG0)
);
// switch matrix multiplexer S1BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S1BEG1 (
    .A0(J2MID_EFb_END0),
    .A1(JE2END0),
    .A2(LF_O),
    .A3(J_l_EF_END2),
    .S0(ConfigBits[338]),
    .S0N(ConfigBits_N[338]),
    .S1(ConfigBits[339]),
    .S1N(ConfigBits_N[339]),
    .X(S1BEG1)
);
// switch matrix multiplexer S1BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S1BEG2 (
    .A0(J2MID_GHb_END1),
    .A1(JE2END1),
    .A2(LG_O),
    .A3(J_l_GH_END3),
    .S0(ConfigBits[340]),
    .S0N(ConfigBits_N[340]),
    .S1(ConfigBits[341]),
    .S1N(ConfigBits_N[341]),
    .X(S1BEG2)
);
// switch matrix multiplexer S1BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S1BEG3 (
    .A0(J2MID_ABb_END2),
    .A1(JE2END2),
    .A2(LH_O),
    .A3(J_l_AB_END0),
    .S0(ConfigBits[342]),
    .S0N(ConfigBits_N[342]),
    .S1(ConfigBits[343]),
    .S1N(ConfigBits_N[343]),
    .X(S1BEG3)
);
// switch matrix multiplexer W1BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_W1BEG0 (
    .A0(J2MID_CDb_END3),
    .A1(JS2END3),
    .A2(LF_O),
    .A3(J_l_CD_END1),
    .S0(ConfigBits[344]),
    .S0N(ConfigBits_N[344]),
    .S1(ConfigBits[345]),
    .S1N(ConfigBits_N[345]),
    .X(W1BEG0)
);
// switch matrix multiplexer W1BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_W1BEG1 (
    .A0(J2MID_EFb_END0),
    .A1(JS2END0),
    .A2(LG_O),
    .A3(J_l_EF_END2),
    .S0(ConfigBits[346]),
    .S0N(ConfigBits_N[346]),
    .S1(ConfigBits[347]),
    .S1N(ConfigBits_N[347]),
    .X(W1BEG1)
);
// switch matrix multiplexer W1BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_W1BEG2 (
    .A0(J2MID_GHb_END1),
    .A1(JS2END1),
    .A2(LH_O),
    .A3(J_l_GH_END3),
    .S0(ConfigBits[348]),
    .S0N(ConfigBits_N[348]),
    .S1(ConfigBits[349]),
    .S1N(ConfigBits_N[349]),
    .X(W1BEG2)
);
// switch matrix multiplexer W1BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_W1BEG3 (
    .A0(J2MID_ABb_END2),
    .A1(JS2END2),
    .A2(LA_O),
    .A3(J_l_AB_END0),
    .S0(ConfigBits[350]),
    .S0N(ConfigBits_N[350]),
    .S1(ConfigBits[351]),
    .S1N(ConfigBits_N[351]),
    .X(W1BEG3)
);
// switch matrix multiplexer N4BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N4BEG0 (
    .A0(LE_O),
    .A1(E6END1),
    .A2(N2END2),
    .A3(N4END1),
    .S0(ConfigBits[352]),
    .S0N(ConfigBits_N[352]),
    .S1(ConfigBits[353]),
    .S1N(ConfigBits_N[353]),
    .X(N4BEG0)
);
// switch matrix multiplexer N4BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N4BEG1 (
    .A0(LF_O),
    .A1(E6END0),
    .A2(N2END3),
    .A3(N4END2),
    .S0(ConfigBits[354]),
    .S0N(ConfigBits_N[354]),
    .S1(ConfigBits[355]),
    .S1N(ConfigBits_N[355]),
    .X(N4BEG1)
);
// switch matrix multiplexer N4BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N4BEG2 (
    .A0(LG_O),
    .A1(W6END1),
    .A2(N2END0),
    .A3(N4END3),
    .S0(ConfigBits[356]),
    .S0N(ConfigBits_N[356]),
    .S1(ConfigBits[357]),
    .S1N(ConfigBits_N[357]),
    .X(N4BEG2)
);
// switch matrix multiplexer N4BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_N4BEG3 (
    .A0(LH_O),
    .A1(W6END0),
    .A2(N2END1),
    .A3(N4END0),
    .S0(ConfigBits[358]),
    .S0N(ConfigBits_N[358]),
    .S1(ConfigBits[359]),
    .S1N(ConfigBits_N[359]),
    .X(N4BEG3)
);
// switch matrix multiplexer S4BEG0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S4BEG0 (
    .A0(LA_O),
    .A1(E6END1),
    .A2(S2END2),
    .A3(S4END1),
    .S0(ConfigBits[360]),
    .S0N(ConfigBits_N[360]),
    .S1(ConfigBits[361]),
    .S1N(ConfigBits_N[361]),
    .X(S4BEG0)
);
// switch matrix multiplexer S4BEG1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S4BEG1 (
    .A0(LB_O),
    .A1(E6END0),
    .A2(S2END3),
    .A3(S4END2),
    .S0(ConfigBits[362]),
    .S0N(ConfigBits_N[362]),
    .S1(ConfigBits[363]),
    .S1N(ConfigBits_N[363]),
    .X(S4BEG1)
);
// switch matrix multiplexer S4BEG2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S4BEG2 (
    .A0(LC_O),
    .A1(W6END1),
    .A2(S2END0),
    .A3(S4END3),
    .S0(ConfigBits[364]),
    .S0N(ConfigBits_N[364]),
    .S1(ConfigBits[365]),
    .S1N(ConfigBits_N[365]),
    .X(S4BEG2)
);
// switch matrix multiplexer S4BEG3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S4BEG3 (
    .A0(LD_O),
    .A1(W6END0),
    .A2(S2END1),
    .A3(S4END0),
    .S0(ConfigBits[366]),
    .S0N(ConfigBits_N[366]),
    .S1(ConfigBits[367]),
    .S1N(ConfigBits_N[367]),
    .X(S4BEG3)
);
// switch matrix multiplexer E6BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_E6BEG0 (
    .A0(M_AH),
    .A1(M_AB),
    .A2(W1END3),
    .A3(E1END3),
    .A4(J2MID_GHb_END1),
    .A5(J2MID_EFb_END1),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[368]),
    .S0N(ConfigBits_N[368]),
    .S1(ConfigBits[369]),
    .S1N(ConfigBits_N[369]),
    .S2(ConfigBits[370]),
    .S2N(ConfigBits_N[370]),
    .S3(ConfigBits[371]),
    .S3N(ConfigBits_N[371]),
    .X(E6BEG0)
);
// switch matrix multiplexer E6BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_E6BEG1 (
    .A0(M_EF),
    .A1(M_AD),
    .A2(W1END2),
    .A3(E1END2),
    .A4(J2MID_GHa_END2),
    .A5(J2MID_EFa_END2),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[372]),
    .S0N(ConfigBits_N[372]),
    .S1(ConfigBits[373]),
    .S1N(ConfigBits_N[373]),
    .S2(ConfigBits[374]),
    .S2N(ConfigBits_N[374]),
    .S3(ConfigBits[375]),
    .S3N(ConfigBits_N[375]),
    .X(E6BEG1)
);
// switch matrix multiplexer W6BEG0 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_W6BEG0 (
    .A0(M_AH),
    .A1(M_AB),
    .A2(W1END3),
    .A3(E1END3),
    .A4(J2MID_GHb_END1),
    .A5(J2MID_EFb_END1),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[376]),
    .S0N(ConfigBits_N[376]),
    .S1(ConfigBits[377]),
    .S1N(ConfigBits_N[377]),
    .S2(ConfigBits[378]),
    .S2N(ConfigBits_N[378]),
    .S3(ConfigBits[379]),
    .S3N(ConfigBits_N[379]),
    .X(W6BEG0)
);
// switch matrix multiplexer W6BEG1 MUX-16cus_mux161_buf_pack #(
    .WIDTH(1)
) inst_cus_mux161_buf_pack_W6BEG1 (
    .A0(M_EF),
    .A1(M_AD),
    .A2(W1END2),
    .A3(E1END2),
    .A4(J2MID_GHa_END2),
    .A5(J2MID_EFa_END2),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .A8(LH_O),
    .A9(LG_O),
    .A10(LF_O),
    .A11(LE_O),
    .A12(LD_O),
    .A13(LC_O),
    .A14(LB_O),
    .A15(LA_O),
    .S0(ConfigBits[380]),
    .S0N(ConfigBits_N[380]),
    .S1(ConfigBits[381]),
    .S1N(ConfigBits_N[381]),
    .S2(ConfigBits[382]),
    .S2N(ConfigBits_N[382]),
    .S3(ConfigBits[383]),
    .S3N(ConfigBits_N[383]),
    .X(W6BEG1)
);
// switch matrix multiplexer EE4BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_EE4BEG0 (
    .A0(E1END2),
    .A1(S1END2),
    .A2(N1END2),
    .A3(J2END_GH_END0),
    .A4(LG_O),
    .A5(LF_O),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .S0(ConfigBits[384]),
    .S0N(ConfigBits_N[384]),
    .S1(ConfigBits[385]),
    .S1N(ConfigBits_N[385]),
    .S2(ConfigBits[386]),
    .S2N(ConfigBits_N[386]),
    .X(EE4BEG0)
);
// switch matrix multiplexer EE4BEG1 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_EE4BEG1 (
    .A0(E1END3),
    .A1(S1END3),
    .A2(N1END3),
    .A3(J2END_EF_END0),
    .A4(LH_O),
    .A5(LA_O),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .S0(ConfigBits[387]),
    .S0N(ConfigBits_N[387]),
    .S1(ConfigBits[388]),
    .S1N(ConfigBits_N[388]),
    .S2(ConfigBits[389]),
    .S2N(ConfigBits_N[389]),
    .X(EE4BEG1)
);
// switch matrix multiplexer EE4BEG2 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_EE4BEG2 (
    .A0(E1END0),
    .A1(S1END0),
    .A2(N1END0),
    .A3(J2END_CD_END0),
    .A4(LC_O),
    .A5(LB_O),
    .A6(J2MID_GHb_END1),
    .A7(J2MID_EFb_END1),
    .S0(ConfigBits[390]),
    .S0N(ConfigBits_N[390]),
    .S1(ConfigBits[391]),
    .S1N(ConfigBits_N[391]),
    .S2(ConfigBits[392]),
    .S2N(ConfigBits_N[392]),
    .X(EE4BEG2)
);
// switch matrix multiplexer EE4BEG3 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_EE4BEG3 (
    .A0(E1END1),
    .A1(S1END1),
    .A2(N1END1),
    .A3(J2END_AB_END0),
    .A4(LE_O),
    .A5(LD_O),
    .A6(J2MID_GHa_END2),
    .A7(J2MID_EFa_END2),
    .S0(ConfigBits[393]),
    .S0N(ConfigBits_N[393]),
    .S1(ConfigBits[394]),
    .S1N(ConfigBits_N[394]),
    .S2(ConfigBits[395]),
    .S2N(ConfigBits_N[395]),
    .X(EE4BEG3)
);
// switch matrix multiplexer WW4BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_WW4BEG0 (
    .A0(W1END2),
    .A1(S1END2),
    .A2(N1END2),
    .A3(J2END_GH_END2),
    .A4(LG_O),
    .A5(LF_O),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .S0(ConfigBits[396]),
    .S0N(ConfigBits_N[396]),
    .S1(ConfigBits[397]),
    .S1N(ConfigBits_N[397]),
    .S2(ConfigBits[398]),
    .S2N(ConfigBits_N[398]),
    .X(WW4BEG0)
);
// switch matrix multiplexer WW4BEG1 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_WW4BEG1 (
    .A0(W1END3),
    .A1(S1END3),
    .A2(N1END3),
    .A3(J2END_EF_END2),
    .A4(LH_O),
    .A5(LA_O),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .S0(ConfigBits[399]),
    .S0N(ConfigBits_N[399]),
    .S1(ConfigBits[400]),
    .S1N(ConfigBits_N[400]),
    .S2(ConfigBits[401]),
    .S2N(ConfigBits_N[401]),
    .X(WW4BEG1)
);
// switch matrix multiplexer WW4BEG2 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_WW4BEG2 (
    .A0(W1END0),
    .A1(S1END0),
    .A2(N1END0),
    .A3(J2END_CD_END2),
    .A4(LC_O),
    .A5(LB_O),
    .A6(J2MID_GHb_END1),
    .A7(J2MID_EFb_END1),
    .S0(ConfigBits[402]),
    .S0N(ConfigBits_N[402]),
    .S1(ConfigBits[403]),
    .S1N(ConfigBits_N[403]),
    .S2(ConfigBits[404]),
    .S2N(ConfigBits_N[404]),
    .X(WW4BEG2)
);
// switch matrix multiplexer WW4BEG3 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_WW4BEG3 (
    .A0(W1END1),
    .A1(S1END1),
    .A2(N1END1),
    .A3(J2END_AB_END2),
    .A4(LE_O),
    .A5(LD_O),
    .A6(J2MID_GHa_END2),
    .A7(J2MID_EFa_END2),
    .S0(ConfigBits[405]),
    .S0N(ConfigBits_N[405]),
    .S1(ConfigBits[406]),
    .S1N(ConfigBits_N[406]),
    .S2(ConfigBits[407]),
    .S2N(ConfigBits_N[407]),
    .X(WW4BEG3)
);
// switch matrix multiplexer NN4BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_NN4BEG0 (
    .A0(N1END2),
    .A1(W1END2),
    .A2(E1END2),
    .A3(J2END_GH_END1),
    .A4(LG_O),
    .A5(LF_O),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .S0(ConfigBits[408]),
    .S0N(ConfigBits_N[408]),
    .S1(ConfigBits[409]),
    .S1N(ConfigBits_N[409]),
    .S2(ConfigBits[410]),
    .S2N(ConfigBits_N[410]),
    .X(NN4BEG0)
);
// switch matrix multiplexer NN4BEG1 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_NN4BEG1 (
    .A0(N1END3),
    .A1(W1END3),
    .A2(E1END3),
    .A3(J2END_EF_END1),
    .A4(LH_O),
    .A5(LA_O),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .S0(ConfigBits[411]),
    .S0N(ConfigBits_N[411]),
    .S1(ConfigBits[412]),
    .S1N(ConfigBits_N[412]),
    .S2(ConfigBits[413]),
    .S2N(ConfigBits_N[413]),
    .X(NN4BEG1)
);
// switch matrix multiplexer NN4BEG2 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_NN4BEG2 (
    .A0(N1END0),
    .A1(W1END0),
    .A2(E1END0),
    .A3(J2END_CD_END1),
    .A4(LC_O),
    .A5(LB_O),
    .A6(J2MID_GHb_END1),
    .A7(J2MID_EFb_END1),
    .S0(ConfigBits[414]),
    .S0N(ConfigBits_N[414]),
    .S1(ConfigBits[415]),
    .S1N(ConfigBits_N[415]),
    .S2(ConfigBits[416]),
    .S2N(ConfigBits_N[416]),
    .X(NN4BEG2)
);
// switch matrix multiplexer NN4BEG3 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_NN4BEG3 (
    .A0(N1END1),
    .A1(W1END1),
    .A2(E1END1),
    .A3(J2END_AB_END1),
    .A4(LE_O),
    .A5(LD_O),
    .A6(J2MID_GHa_END2),
    .A7(J2MID_EFa_END2),
    .S0(ConfigBits[417]),
    .S0N(ConfigBits_N[417]),
    .S1(ConfigBits[418]),
    .S1N(ConfigBits_N[418]),
    .S2(ConfigBits[419]),
    .S2N(ConfigBits_N[419]),
    .X(NN4BEG3)
);
// switch matrix multiplexer SS4BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_SS4BEG0 (
    .A0(N1END2),
    .A1(W1END2),
    .A2(E1END2),
    .A3(J2END_GH_END3),
    .A4(LG_O),
    .A5(LF_O),
    .A6(J2MID_CDb_END1),
    .A7(J2MID_ABb_END1),
    .S0(ConfigBits[420]),
    .S0N(ConfigBits_N[420]),
    .S1(ConfigBits[421]),
    .S1N(ConfigBits_N[421]),
    .S2(ConfigBits[422]),
    .S2N(ConfigBits_N[422]),
    .X(SS4BEG0)
);
// switch matrix multiplexer SS4BEG1 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_SS4BEG1 (
    .A0(N1END3),
    .A1(W1END3),
    .A2(E1END3),
    .A3(J2END_EF_END3),
    .A4(LH_O),
    .A5(LA_O),
    .A6(J2MID_CDa_END2),
    .A7(J2MID_ABa_END2),
    .S0(ConfigBits[423]),
    .S0N(ConfigBits_N[423]),
    .S1(ConfigBits[424]),
    .S1N(ConfigBits_N[424]),
    .S2(ConfigBits[425]),
    .S2N(ConfigBits_N[425]),
    .X(SS4BEG1)
);
// switch matrix multiplexer SS4BEG2 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_SS4BEG2 (
    .A0(N1END0),
    .A1(W1END0),
    .A2(E1END0),
    .A3(J2END_CD_END3),
    .A4(LC_O),
    .A5(LB_O),
    .A6(J2MID_GHb_END1),
    .A7(J2MID_EFb_END1),
    .S0(ConfigBits[426]),
    .S0N(ConfigBits_N[426]),
    .S1(ConfigBits[427]),
    .S1N(ConfigBits_N[427]),
    .S2(ConfigBits[428]),
    .S2N(ConfigBits_N[428]),
    .X(SS4BEG2)
);
// switch matrix multiplexer SS4BEG3 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_SS4BEG3 (
    .A0(N1END1),
    .A1(W1END1),
    .A2(E1END1),
    .A3(J2END_AB_END3),
    .A4(LE_O),
    .A5(LD_O),
    .A6(J2MID_GHa_END2),
    .A7(J2MID_EFa_END2),
    .S0(ConfigBits[429]),
    .S0N(ConfigBits_N[429]),
    .S1(ConfigBits[430]),
    .S1N(ConfigBits_N[430]),
    .S2(ConfigBits[431]),
    .S2N(ConfigBits_N[431]),
    .X(SS4BEG3)
);
// switch matrix multiplexer A MUX-1assign A = LA_O;// switch matrix multiplexer B MUX-1assign B = LB_O;// switch matrix multiplexer C MUX-1assign C = LC_O;// switch matrix multiplexer D MUX-1assign D = LD_O;// switch matrix multiplexer E MUX-1assign E = LE_O;// switch matrix multiplexer F MUX-1assign F = LF_O;// switch matrix multiplexer G MUX-1assign G = LG_O;// switch matrix multiplexer H MUX-1assign H = LH_O;// switch matrix multiplexer S0 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S0 (
    .A0(JW2END4),
    .A1(JS2END4),
    .A2(JE2END4),
    .A3(JN2END4),
    .S0(ConfigBits[432]),
    .S0N(ConfigBits_N[432]),
    .S1(ConfigBits[433]),
    .S1N(ConfigBits_N[433]),
    .X(S0)
);
// switch matrix multiplexer S1 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S1 (
    .A0(JW2END5),
    .A1(JS2END5),
    .A2(JE2END5),
    .A3(JN2END5),
    .S0(ConfigBits[434]),
    .S0N(ConfigBits_N[434]),
    .S1(ConfigBits[435]),
    .S1N(ConfigBits_N[435]),
    .X(S1)
);
// switch matrix multiplexer S2 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S2 (
    .A0(JW2END6),
    .A1(JS2END6),
    .A2(JE2END6),
    .A3(JN2END6),
    .S0(ConfigBits[436]),
    .S0N(ConfigBits_N[436]),
    .S1(ConfigBits[437]),
    .S1N(ConfigBits_N[437]),
    .X(S2)
);
// switch matrix multiplexer S3 MUX-4cus_mux41_buf_pack #(
    .WIDTH(1)
) inst_cus_mux41_buf_pack_S3 (
    .A0(JW2END7),
    .A1(JS2END7),
    .A2(JE2END7),
    .A3(JN2END7),
    .S0(ConfigBits[438]),
    .S0N(ConfigBits_N[438]),
    .S1(ConfigBits[439]),
    .S1N(ConfigBits_N[439]),
    .X(S3)
);
// switch matrix multiplexer LA_Ci MUX-1assign LA_Ci = Ci0;// switch matrix multiplexer LB_Ci MUX-1assign LB_Ci = LA_Co;// switch matrix multiplexer LC_Ci MUX-1assign LC_Ci = LB_Co;// switch matrix multiplexer LD_Ci MUX-1assign LD_Ci = LC_Co;// switch matrix multiplexer LE_Ci MUX-1assign LE_Ci = LD_Co;// switch matrix multiplexer LF_Ci MUX-1assign LF_Ci = LE_Co;// switch matrix multiplexer LG_Ci MUX-1assign LG_Ci = LF_Co;// switch matrix multiplexer LH_Ci MUX-1assign LH_Ci = LG_Co;// switch matrix multiplexer Co0 MUX-1assign Co0 = LH_Co;// switch matrix multiplexer J_SR_BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_J_SR_BEG0 (
    .A0(JW2END1),
    .A1(JS2END1),
    .A2(JE2END1),
    .A3(JN2END1),
    .A4(J2MID_GHa_END0),
    .A5(J2MID_EFb_END0),
    .A6(J2MID_CDb_END0),
    .A7(J2MID_ABb_END0),
    .S0(ConfigBits[440]),
    .S0N(ConfigBits_N[440]),
    .S1(ConfigBits[441]),
    .S1N(ConfigBits_N[441]),
    .S2(ConfigBits[442]),
    .S2N(ConfigBits_N[442]),
    .X(J_SR_BEG0)
);
// switch matrix multiplexer J_EN_BEG0 MUX-8cus_mux81_buf_pack #(
    .WIDTH(1)
) inst_cus_mux81_buf_pack_J_EN_BEG0 (
    .A0(JW2END2),
    .A1(JS2END2),
    .A2(JE2END2),
    .A3(JN2END2),
    .A4(J2MID_GHa_END3),
    .A5(J2MID_EFb_END3),
    .A6(J2MID_CDb_END3),
    .A7(J2MID_ABb_END3),
    .S0(ConfigBits[443]),
    .S0N(ConfigBits_N[443]),
    .S1(ConfigBits[444]),
    .S1N(ConfigBits_N[444]),
    .S2(ConfigBits[445]),
    .S2N(ConfigBits_N[445]),
    .X(J_EN_BEG0)
);
// switch matrix multiplexer LA_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LA_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[446]),
    .X(LA_SR)
);
// switch matrix multiplexer LB_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LB_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[447]),
    .X(LB_SR)
);
// switch matrix multiplexer LC_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LC_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[448]),
    .X(LC_SR)
);
// switch matrix multiplexer LD_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LD_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[449]),
    .X(LD_SR)
);
// switch matrix multiplexer LE_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LE_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[450]),
    .X(LE_SR)
);
// switch matrix multiplexer LF_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LF_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[451]),
    .X(LF_SR)
);
// switch matrix multiplexer LG_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LG_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[452]),
    .X(LG_SR)
);
// switch matrix multiplexer LH_SR MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LH_SR (
    .A0(GND0),
    .A1(J_SR_END0),
    .S(ConfigBits[453]),
    .X(LH_SR)
);
// switch matrix multiplexer LA_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LA_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[454]),
    .X(LA_EN)
);
// switch matrix multiplexer LB_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LB_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[455]),
    .X(LB_EN)
);
// switch matrix multiplexer LC_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LC_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[456]),
    .X(LC_EN)
);
// switch matrix multiplexer LD_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LD_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[457]),
    .X(LD_EN)
);
// switch matrix multiplexer LE_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LE_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[458]),
    .X(LE_EN)
);
// switch matrix multiplexer LF_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LF_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[459]),
    .X(LF_EN)
);
// switch matrix multiplexer LG_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LG_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[460]),
    .X(LG_EN)
);
// switch matrix multiplexer LH_EN MUX-2cus_mux21_pack #(
    .WIDTH(1)
) inst_cus_mux21_pack_LH_EN (
    .A0(VCC0),
    .A1(J_EN_END0),
    .S(ConfigBits[461]),
    .X(LH_EN)
);

endmodule
