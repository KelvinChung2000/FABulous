module cap #(parameter WIDTH=32);

localparam add_op = 0;
localparam ashr_op = 1;
localparam const_op = 2;
localparam icmp_op = 3;
localparam io_width_1_op = 4;
localparam mul_op = 5;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const1;
wire[WIDTH-1:0] i2_mul1;
wire[WIDTH-1:0] i2_add1;
wire[WIDTH-1:0] i3_load;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i4_mul;
wire[WIDTH-1:0] c1;
wire[WIDTH-1:0] i5_load;
wire[WIDTH-1:0] i6_mul;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i7_ashr;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i8_data_size1;
wire[WIDTH-1:0] i8_mul1;
wire[WIDTH-1:0] i8_add1;
wire[WIDTH-1:0] i9_load;
wire[WIDTH-1:0] i10_mul;
wire[WIDTH-1:0] i11_ashr;
wire[WIDTH-1:0] i12_mul;
wire[WIDTH-1:0] i13_mul;
wire[WIDTH-1:0] i14_mul;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i15_data_size1;
wire[WIDTH-1:0] i15_mul1;
wire[WIDTH-1:0] i15_add1;
wire[WIDTH-1:0] const6;
wire[WIDTH-1:0] i17_add;
wire[WIDTH-1:0] input0;
wire i18_icmp;
wire[WIDTH-1:0] const3_dup_1;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const1_alu;
wire[WIDTH-1:0] i2_mul1_alu;
wire[WIDTH-1:0] i2_add1_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i4_mul_alu;
wire[WIDTH-1:0] i6_mul_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i7_ashr_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i8_data_size1_alu;
wire[WIDTH-1:0] i8_mul1_alu;
wire[WIDTH-1:0] i8_add1_alu;
wire[WIDTH-1:0] i10_mul_alu;
wire[WIDTH-1:0] i11_ashr_alu;
wire[WIDTH-1:0] i12_mul_alu;
wire[WIDTH-1:0] i13_mul_alu;
wire[WIDTH-1:0] i14_mul_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i15_data_size1_alu;
wire[WIDTH-1:0] i15_mul1_alu;
wire[WIDTH-1:0] i15_add1_alu;
wire[WIDTH-1:0] const6_alu;
wire[WIDTH-1:0] i17_add_alu;
wire[WIDTH-1:0] const3_dup_1_alu;
wire[WIDTH-1:0] i16_store;
wire[WIDTH-1:0] i19_br;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(8)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const1(.const_out(const1));
ALU #(.ALU_func(mul_op)) inst_i2_mul1(.data_in1(const0), .data_in2(i17_add), .data_in3(), .data_out(i2_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i2_mul1_reg(.reg_in(i2_mul1_alu), .reg_out(i2_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i2_add1(.data_in1(const1), .data_in2(i2_mul1), .data_in3(), .data_out(i2_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i2_add1_reg(.reg_in(i2_add1_alu), .reg_out(i2_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i3_load(.addr0(i2_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i3_load));
const_unit #(.ConfigBits(3)) inst_const2(.const_out(const2));
ALU #(.ALU_func(mul_op)) inst_i4_mul(.data_in1(i3_load), .data_in2(const2), .data_in3(), .data_out(i4_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_mul_reg(.reg_in(i4_mul_alu), .reg_out(i4_mul), .en(global_en), .rst(global_rst));
(* keep *) IO inst_c1(.from_fabric(), .in(), .to_fabric(c1), .out());
(* keep *)Mem #(.config_bits(0)) inst_i5_load(.addr0(c1), .reset(global_rst), .write_data(), .write_en(), .read_data(i5_load));
ALU #(.ALU_func(mul_op)) inst_i6_mul(.data_in1(i4_mul), .data_in2(i5_load), .data_in3(), .data_out(i6_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_mul_reg(.reg_in(i6_mul_alu), .reg_out(i6_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2)) inst_const3(.const_out(const3));
ALU #(.ALU_func(ashr_op)) inst_i7_ashr(.data_in1(i6_mul), .data_in2(const3), .data_in3(), .data_out(i7_ashr_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_ashr_reg(.reg_in(i7_ashr_alu), .reg_out(i7_ashr), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(3584)) inst_const4(.const_out(const4));
const_unit #(.ConfigBits(4)) inst_i8_data_size1(.const_out(i8_data_size1));
ALU #(.ALU_func(mul_op)) inst_i8_mul1(.data_in1(i8_data_size1), .data_in2(i17_add), .data_in3(), .data_out(i8_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_mul1_reg(.reg_in(i8_mul1_alu), .reg_out(i8_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i8_add1(.data_in1(const4), .data_in2(i8_mul1), .data_in3(), .data_out(i8_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_add1_reg(.reg_in(i8_add1_alu), .reg_out(i8_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i9_load(.addr0(i8_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i9_load));
ALU #(.ALU_func(mul_op)) inst_i10_mul(.data_in1(i4_mul), .data_in2(i9_load), .data_in3(), .data_out(i10_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_mul_reg(.reg_in(i10_mul_alu), .reg_out(i10_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(ashr_op)) inst_i11_ashr(.data_in1(i10_mul), .data_in2(const3_dup_1), .data_in3(), .data_out(i11_ashr_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_ashr_reg(.reg_in(i11_ashr_alu), .reg_out(i11_ashr), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i12_mul(.data_in1(i3_load), .data_in2(i5_load), .data_in3(), .data_out(i12_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_mul_reg(.reg_in(i12_mul_alu), .reg_out(i12_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i13_mul(.data_in1(i7_ashr), .data_in2(i12_mul), .data_in3(), .data_out(i13_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i13_mul_reg(.reg_in(i13_mul_alu), .reg_out(i13_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i14_mul(.data_in1(i11_ashr), .data_in2(i13_mul), .data_in3(), .data_out(i14_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_mul_reg(.reg_in(i14_mul_alu), .reg_out(i14_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2816)) inst_const5(.const_out(const5));
const_unit #(.ConfigBits(4)) inst_i15_data_size1(.const_out(i15_data_size1));
ALU #(.ALU_func(mul_op)) inst_i15_mul1(.data_in1(i15_data_size1), .data_in2(i17_add), .data_in3(), .data_out(i15_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_mul1_reg(.reg_in(i15_mul1_alu), .reg_out(i15_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i15_add1(.data_in1(const5), .data_in2(i15_mul1), .data_in3(), .data_out(i15_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_add1_reg(.reg_in(i15_add1_alu), .reg_out(i15_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i16_store(.addr0(i14_mul), .reset(global_rst), .write_data(i15_add1), .write_en(), .read_data(i16_store));
const_unit #(.ConfigBits(1)) inst_const6(.const_out(const6));
ALU #(.ALU_func(add_op)) inst_i17_add(.data_in1(const6), .data_in2(i17_add), .data_in3(), .data_out(i17_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i17_add_reg(.reg_in(i17_add_alu), .reg_out(i17_add), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i18_icmp(.A(i17_add), .B(input0), .Y(i18_icmp));
(* keep *) IO_WIDTH_1 inst_i19_br(.from_fabric(i18_icmp), .in(), .to_fabric(), .out());
const_unit #(.ConfigBits(2)) inst_const3_dup_1(.const_out(const3_dup_1));

endmodule
