module ALU #(
    parameter NoConfigBits = 3,
    parameter WIDTH = 32
) (
    input wire rst,
    input wire en,
    (* FABulous, USER_CLK *) input wire clk,
    (* FABulous, BUS *) input wire [WIDTH-1:0] data_in1,
    (* FABulous, BUS *) input wire [WIDTH-1:0] data_in2,
    (* FABulous, BUS *) input wire [WIDTH-1:0] data_in3,
    (* FABulous, BUS *) output reg [WIDTH-1:0] data_out,
    (* FABulous, CONFIG_BIT, FEATURE="ALU", FEATURE_MAP="std_add(left=>data_in1, right=>data_in2, out=>data_out);" *) input [NoConfigBits:0] ConfigBits
);
  // Define operation codes
  localparam ADD = 3'b000;
  localparam SUB = 3'b001;
  localparam AND = 3'b010;
  localparam OR = 3'b011;
  localparam XOR = 3'b100;
  localparam MUL = 3'b101;

  always @(*) begin
    if (rst) begin
      data_out = 8'b0;
    end else if (en) begin
      case (ConfigBits)
        ADD: data_out = data_in1 + data_in2;
        SUB: data_out = data_in1 - data_in2;
        AND: data_out = data_in1 & data_in2;
        OR: data_out = data_in1 | data_in2;
        XOR: data_out = data_in1 ^ data_in2;
        MUL: data_out = data_in1 * data_in2;
        default: data_out = 8'b0;
      endcase
    end
  end


endmodule
