(* blackbox *)
module IO #(

)(
    input [31:0] from_fabric,
    input [31:0] in,
    output [31:0] to_fabric,
    output [31:0] out
);

endmodule
