(* blackbox *)
module const_unit #(
    parameter ConfigBits = 0
)(
    output [31:0] const_out
);

endmodule

