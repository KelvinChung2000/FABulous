module simple2 #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] a;
wire[WIDTH-1:0] i2_load;
wire[WIDTH-1:0] i3_data_size1;
wire[WIDTH-1:0] i3_mul1;
wire[WIDTH-1:0] i3_add1;
wire[WIDTH-1:0] i4_load;
wire[WIDTH-1:0] b;
wire[WIDTH-1:0] i5_load;
wire[WIDTH-1:0] i6_data_size1;
wire[WIDTH-1:0] i6_mul1;
wire[WIDTH-1:0] i6_add1;
wire[WIDTH-1:0] i7_load;
wire[WIDTH-1:0] i8_mul;
wire[WIDTH-1:0] input0;
wire[WIDTH-1:0] i9_data_size1;
wire[WIDTH-1:0] i9_mul1;
wire[WIDTH-1:0] i9_add1;
wire[WIDTH-1:0] i9_data_size2;
wire[WIDTH-1:0] i9_mul2;
wire[WIDTH-1:0] i9_add2;
wire[WIDTH-1:0] const1;
wire[WIDTH-1:0] i11_add;
wire[WIDTH-1:0] const2;
wire i12_icmp;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] i3_data_size1_alu;
wire[WIDTH-1:0] i3_mul1_alu;
wire[WIDTH-1:0] i3_add1_alu;
wire[WIDTH-1:0] i6_data_size1_alu;
wire[WIDTH-1:0] i6_mul1_alu;
wire[WIDTH-1:0] i6_add1_alu;
wire[WIDTH-1:0] i8_mul_alu;
wire[WIDTH-1:0] i9_data_size1_alu;
wire[WIDTH-1:0] i9_mul1_alu;
wire[WIDTH-1:0] i9_add1_alu;
wire[WIDTH-1:0] i9_data_size2_alu;
wire[WIDTH-1:0] i9_mul2_alu;
wire[WIDTH-1:0] i9_add2_alu;
wire[WIDTH-1:0] const1_alu;
wire[WIDTH-1:0] i11_add_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i10_store;
wire[WIDTH-1:0] i13_br;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(0)) inst_const0(.const_out(const0));
(* keep *) IO inst_a(.from_fabric(), .in(), .to_fabric(a), .out());
(* keep *)Mem #(.config_bits(0)) inst_i2_load(.addr0(a), .reset(global_rst), .write_data(), .write_en(), .read_data(i2_load));
const_unit #(.ConfigBits(4)) inst_i3_data_size1(.const_out(i3_data_size1));
ALU #(.ALU_func(mul_op)) inst_i3_mul1(.data_in1(i3_data_size1), .data_in2(i11_add), .data_in3(), .data_out(i3_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_mul1_reg(.reg_in(i3_mul1_alu), .reg_out(i3_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i3_add1(.data_in1(i2_load), .data_in2(i3_mul1), .data_in3(), .data_out(i3_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add1_reg(.reg_in(i3_add1_alu), .reg_out(i3_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i4_load(.addr0(i3_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i4_load));
(* keep *) IO inst_b(.from_fabric(), .in(), .to_fabric(b), .out());
(* keep *)Mem #(.config_bits(0)) inst_i5_load(.addr0(b), .reset(global_rst), .write_data(), .write_en(), .read_data(i5_load));
const_unit #(.ConfigBits(4)) inst_i6_data_size1(.const_out(i6_data_size1));
ALU #(.ALU_func(mul_op)) inst_i6_mul1(.data_in1(i6_data_size1), .data_in2(i11_add), .data_in3(), .data_out(i6_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_mul1_reg(.reg_in(i6_mul1_alu), .reg_out(i6_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i6_add1(.data_in1(i5_load), .data_in2(i6_mul1), .data_in3(), .data_out(i6_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add1_reg(.reg_in(i6_add1_alu), .reg_out(i6_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i7_load(.addr0(i6_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i7_load));
ALU #(.ALU_func(mul_op)) inst_i8_mul(.data_in1(i4_load), .data_in2(i7_load), .data_in3(), .data_out(i8_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_mul_reg(.reg_in(i8_mul_alu), .reg_out(i8_mul), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
const_unit #(.ConfigBits(80)) inst_i9_data_size1(.const_out(i9_data_size1));
ALU #(.ALU_func(mul_op)) inst_i9_mul1(.data_in1(const0), .data_in2(i9_data_size1), .data_in3(), .data_out(i9_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_mul1_reg(.reg_in(i9_mul1_alu), .reg_out(i9_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i9_add1(.data_in1(input0), .data_in2(i9_mul1), .data_in3(), .data_out(i9_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add1_reg(.reg_in(i9_add1_alu), .reg_out(i9_add1), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i9_data_size2(.const_out(i9_data_size2));
ALU #(.ALU_func(mul_op)) inst_i9_mul2(.data_in1(i9_data_size2), .data_in2(i11_add), .data_in3(), .data_out(i9_mul2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_mul2_reg(.reg_in(i9_mul2_alu), .reg_out(i9_mul2), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i9_add2(.data_in1(i9_add1), .data_in2(i9_mul2), .data_in3(), .data_out(i9_add2_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add2_reg(.reg_in(i9_add2_alu), .reg_out(i9_add2), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i10_store(.addr0(i8_mul), .reset(global_rst), .write_data(i9_add2), .write_en(), .read_data(i10_store));
const_unit #(.ConfigBits(1)) inst_const1(.const_out(const1));
ALU #(.ALU_func(add_op)) inst_i11_add(.data_in1(const1), .data_in2(i11_add), .data_in3(), .data_out(i11_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_add_reg(.reg_in(i11_add_alu), .reg_out(i11_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(20)) inst_const2(.const_out(const2));
compare #(.conf(0)) inst_i12_icmp(.A(i11_add), .B(const2), .Y(i12_icmp));
(* keep *) IO_WIDTH_1 inst_i13_br(.from_fabric(i12_icmp), .in(), .to_fabric(), .out());

endmodule
