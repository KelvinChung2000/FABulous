module eFPGA_top
    #(
        parameter include_eFPGA=1,
        parameter NumberOfRows=14,
        parameter NumberOfCols=10,
        parameter FrameBitsPerRow=32,
        parameter MaxFramesPerCol=20,
        parameter desync_flag=20,
        parameter FrameSelectWidth=5,
        parameter RowSelectWidth=5
    )
    (
        //External IO port
        output [55:0] A_config_C,
        output [55:0] B_config_C,
        output [55:0] Config_accessC,
        output [27:0] I_top,
        input [27:0] O_top,
        output [27:0] T_top,
        //Config related ports
        input CLK,
        input resetn,
        input SelfWriteStrobe,
        input [31:0] SelfWriteData,
        input Rx,
        output ComActive,
        output ReceiveLED,
        input s_clk,
        input s_data
);
 //BlockRAM ports

wire[224-1:0] RAM2FAB_D_I;
wire[224-1:0] FAB2RAM_D_O;
wire[112-1:0] FAB2RAM_A_O;
wire[56-1:0] FAB2RAM_C_O;

 //Signal declarations
wire[(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;
wire[(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;
wire[(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;
wire[FrameBitsPerRow-1:0] FrameAddressRegister;
wire LongFrameStrobe;
wire[31:0] LocalWriteData;
wire LocalWriteStrobe;
wire[RowSelectWidth-1:0] RowSelect;
`ifndef EMULATION

eFPGA_Config
    #(
    .RowSelectWidth(RowSelectWidth),
    .NumberOfRows(NumberOfRows),
    .desync_flag(desync_flag),
    .FrameBitsPerRow(FrameBitsPerRow)
    )
    eFPGA_Config_inst
    (
    .CLK(CLK),
    .resetn(resetn),
    .Rx(Rx),
    .ComActive(ComActive),
    .ReceiveLED(ReceiveLED),
    .s_clk(s_clk),
    .s_data(s_data),
    .SelfWriteData(SelfWriteData),
    .SelfWriteStrobe(SelfWriteStrobe),
    .ConfigWriteData(LocalWriteData),
    .ConfigWriteStrobe(LocalWriteStrobe),
    .FrameAddressRegister(FrameAddressRegister),
    .LongFrameStrobe(LongFrameStrobe),
    .RowSelect(RowSelect)
);


Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(1)
    )
    inst_Frame_Data_Reg_0
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[0*FrameBitsPerRow+FrameBitsPerRow-1:0*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(2)
    )
    inst_Frame_Data_Reg_1
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[1*FrameBitsPerRow+FrameBitsPerRow-1:1*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(3)
    )
    inst_Frame_Data_Reg_2
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[2*FrameBitsPerRow+FrameBitsPerRow-1:2*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(4)
    )
    inst_Frame_Data_Reg_3
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[3*FrameBitsPerRow+FrameBitsPerRow-1:3*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(5)
    )
    inst_Frame_Data_Reg_4
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[4*FrameBitsPerRow+FrameBitsPerRow-1:4*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(6)
    )
    inst_Frame_Data_Reg_5
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[5*FrameBitsPerRow+FrameBitsPerRow-1:5*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(7)
    )
    inst_Frame_Data_Reg_6
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[6*FrameBitsPerRow+FrameBitsPerRow-1:6*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(8)
    )
    inst_Frame_Data_Reg_7
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[7*FrameBitsPerRow+FrameBitsPerRow-1:7*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(9)
    )
    inst_Frame_Data_Reg_8
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[8*FrameBitsPerRow+FrameBitsPerRow-1:8*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(10)
    )
    inst_Frame_Data_Reg_9
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[9*FrameBitsPerRow+FrameBitsPerRow-1:9*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(11)
    )
    inst_Frame_Data_Reg_10
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[10*FrameBitsPerRow+FrameBitsPerRow-1:10*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(12)
    )
    inst_Frame_Data_Reg_11
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[11*FrameBitsPerRow+FrameBitsPerRow-1:11*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(13)
    )
    inst_Frame_Data_Reg_12
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[12*FrameBitsPerRow+FrameBitsPerRow-1:12*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(14)
    )
    inst_Frame_Data_Reg_13
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[13*FrameBitsPerRow+FrameBitsPerRow-1:13*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);


Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(0)
    )
    inst_Frame_Select_0
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[0*MaxFramesPerCol+MaxFramesPerCol-1:0*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(1)
    )
    inst_Frame_Select_1
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[1*MaxFramesPerCol+MaxFramesPerCol-1:1*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(2)
    )
    inst_Frame_Select_2
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[2*MaxFramesPerCol+MaxFramesPerCol-1:2*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(3)
    )
    inst_Frame_Select_3
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[3*MaxFramesPerCol+MaxFramesPerCol-1:3*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(4)
    )
    inst_Frame_Select_4
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[4*MaxFramesPerCol+MaxFramesPerCol-1:4*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(5)
    )
    inst_Frame_Select_5
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[5*MaxFramesPerCol+MaxFramesPerCol-1:5*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(6)
    )
    inst_Frame_Select_6
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[6*MaxFramesPerCol+MaxFramesPerCol-1:6*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(7)
    )
    inst_Frame_Select_7
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[7*MaxFramesPerCol+MaxFramesPerCol-1:7*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(8)
    )
    inst_Frame_Select_8
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[8*MaxFramesPerCol+MaxFramesPerCol-1:8*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(9)
    )
    inst_Frame_Select_9
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[9*MaxFramesPerCol+MaxFramesPerCol-1:9*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);


`endif
eFPGA eFPGA_inst (
    .Tile_X0Y14_A_config_C_bit0(A_config_C[0]),
    .Tile_X0Y14_A_config_C_bit1(A_config_C[1]),
    .Tile_X0Y14_A_config_C_bit2(A_config_C[2]),
    .Tile_X0Y14_A_config_C_bit3(A_config_C[3]),
    .Tile_X0Y13_A_config_C_bit0(A_config_C[4]),
    .Tile_X0Y13_A_config_C_bit1(A_config_C[5]),
    .Tile_X0Y13_A_config_C_bit2(A_config_C[6]),
    .Tile_X0Y13_A_config_C_bit3(A_config_C[7]),
    .Tile_X0Y12_A_config_C_bit0(A_config_C[8]),
    .Tile_X0Y12_A_config_C_bit1(A_config_C[9]),
    .Tile_X0Y12_A_config_C_bit2(A_config_C[10]),
    .Tile_X0Y12_A_config_C_bit3(A_config_C[11]),
    .Tile_X0Y11_A_config_C_bit0(A_config_C[12]),
    .Tile_X0Y11_A_config_C_bit1(A_config_C[13]),
    .Tile_X0Y11_A_config_C_bit2(A_config_C[14]),
    .Tile_X0Y11_A_config_C_bit3(A_config_C[15]),
    .Tile_X0Y10_A_config_C_bit0(A_config_C[16]),
    .Tile_X0Y10_A_config_C_bit1(A_config_C[17]),
    .Tile_X0Y10_A_config_C_bit2(A_config_C[18]),
    .Tile_X0Y10_A_config_C_bit3(A_config_C[19]),
    .Tile_X0Y9_A_config_C_bit0(A_config_C[20]),
    .Tile_X0Y9_A_config_C_bit1(A_config_C[21]),
    .Tile_X0Y9_A_config_C_bit2(A_config_C[22]),
    .Tile_X0Y9_A_config_C_bit3(A_config_C[23]),
    .Tile_X0Y8_A_config_C_bit0(A_config_C[24]),
    .Tile_X0Y8_A_config_C_bit1(A_config_C[25]),
    .Tile_X0Y8_A_config_C_bit2(A_config_C[26]),
    .Tile_X0Y8_A_config_C_bit3(A_config_C[27]),
    .Tile_X0Y7_A_config_C_bit0(A_config_C[28]),
    .Tile_X0Y7_A_config_C_bit1(A_config_C[29]),
    .Tile_X0Y7_A_config_C_bit2(A_config_C[30]),
    .Tile_X0Y7_A_config_C_bit3(A_config_C[31]),
    .Tile_X0Y6_A_config_C_bit0(A_config_C[32]),
    .Tile_X0Y6_A_config_C_bit1(A_config_C[33]),
    .Tile_X0Y6_A_config_C_bit2(A_config_C[34]),
    .Tile_X0Y6_A_config_C_bit3(A_config_C[35]),
    .Tile_X0Y5_A_config_C_bit0(A_config_C[36]),
    .Tile_X0Y5_A_config_C_bit1(A_config_C[37]),
    .Tile_X0Y5_A_config_C_bit2(A_config_C[38]),
    .Tile_X0Y5_A_config_C_bit3(A_config_C[39]),
    .Tile_X0Y4_A_config_C_bit0(A_config_C[40]),
    .Tile_X0Y4_A_config_C_bit1(A_config_C[41]),
    .Tile_X0Y4_A_config_C_bit2(A_config_C[42]),
    .Tile_X0Y4_A_config_C_bit3(A_config_C[43]),
    .Tile_X0Y3_A_config_C_bit0(A_config_C[44]),
    .Tile_X0Y3_A_config_C_bit1(A_config_C[45]),
    .Tile_X0Y3_A_config_C_bit2(A_config_C[46]),
    .Tile_X0Y3_A_config_C_bit3(A_config_C[47]),
    .Tile_X0Y2_A_config_C_bit0(A_config_C[48]),
    .Tile_X0Y2_A_config_C_bit1(A_config_C[49]),
    .Tile_X0Y2_A_config_C_bit2(A_config_C[50]),
    .Tile_X0Y2_A_config_C_bit3(A_config_C[51]),
    .Tile_X0Y1_A_config_C_bit0(A_config_C[52]),
    .Tile_X0Y1_A_config_C_bit1(A_config_C[53]),
    .Tile_X0Y1_A_config_C_bit2(A_config_C[54]),
    .Tile_X0Y1_A_config_C_bit3(A_config_C[55]),
    .Tile_X0Y14_B_config_C_bit0(B_config_C[0]),
    .Tile_X0Y14_B_config_C_bit1(B_config_C[1]),
    .Tile_X0Y14_B_config_C_bit2(B_config_C[2]),
    .Tile_X0Y14_B_config_C_bit3(B_config_C[3]),
    .Tile_X0Y13_B_config_C_bit0(B_config_C[4]),
    .Tile_X0Y13_B_config_C_bit1(B_config_C[5]),
    .Tile_X0Y13_B_config_C_bit2(B_config_C[6]),
    .Tile_X0Y13_B_config_C_bit3(B_config_C[7]),
    .Tile_X0Y12_B_config_C_bit0(B_config_C[8]),
    .Tile_X0Y12_B_config_C_bit1(B_config_C[9]),
    .Tile_X0Y12_B_config_C_bit2(B_config_C[10]),
    .Tile_X0Y12_B_config_C_bit3(B_config_C[11]),
    .Tile_X0Y11_B_config_C_bit0(B_config_C[12]),
    .Tile_X0Y11_B_config_C_bit1(B_config_C[13]),
    .Tile_X0Y11_B_config_C_bit2(B_config_C[14]),
    .Tile_X0Y11_B_config_C_bit3(B_config_C[15]),
    .Tile_X0Y10_B_config_C_bit0(B_config_C[16]),
    .Tile_X0Y10_B_config_C_bit1(B_config_C[17]),
    .Tile_X0Y10_B_config_C_bit2(B_config_C[18]),
    .Tile_X0Y10_B_config_C_bit3(B_config_C[19]),
    .Tile_X0Y9_B_config_C_bit0(B_config_C[20]),
    .Tile_X0Y9_B_config_C_bit1(B_config_C[21]),
    .Tile_X0Y9_B_config_C_bit2(B_config_C[22]),
    .Tile_X0Y9_B_config_C_bit3(B_config_C[23]),
    .Tile_X0Y8_B_config_C_bit0(B_config_C[24]),
    .Tile_X0Y8_B_config_C_bit1(B_config_C[25]),
    .Tile_X0Y8_B_config_C_bit2(B_config_C[26]),
    .Tile_X0Y8_B_config_C_bit3(B_config_C[27]),
    .Tile_X0Y7_B_config_C_bit0(B_config_C[28]),
    .Tile_X0Y7_B_config_C_bit1(B_config_C[29]),
    .Tile_X0Y7_B_config_C_bit2(B_config_C[30]),
    .Tile_X0Y7_B_config_C_bit3(B_config_C[31]),
    .Tile_X0Y6_B_config_C_bit0(B_config_C[32]),
    .Tile_X0Y6_B_config_C_bit1(B_config_C[33]),
    .Tile_X0Y6_B_config_C_bit2(B_config_C[34]),
    .Tile_X0Y6_B_config_C_bit3(B_config_C[35]),
    .Tile_X0Y5_B_config_C_bit0(B_config_C[36]),
    .Tile_X0Y5_B_config_C_bit1(B_config_C[37]),
    .Tile_X0Y5_B_config_C_bit2(B_config_C[38]),
    .Tile_X0Y5_B_config_C_bit3(B_config_C[39]),
    .Tile_X0Y4_B_config_C_bit0(B_config_C[40]),
    .Tile_X0Y4_B_config_C_bit1(B_config_C[41]),
    .Tile_X0Y4_B_config_C_bit2(B_config_C[42]),
    .Tile_X0Y4_B_config_C_bit3(B_config_C[43]),
    .Tile_X0Y3_B_config_C_bit0(B_config_C[44]),
    .Tile_X0Y3_B_config_C_bit1(B_config_C[45]),
    .Tile_X0Y3_B_config_C_bit2(B_config_C[46]),
    .Tile_X0Y3_B_config_C_bit3(B_config_C[47]),
    .Tile_X0Y2_B_config_C_bit0(B_config_C[48]),
    .Tile_X0Y2_B_config_C_bit1(B_config_C[49]),
    .Tile_X0Y2_B_config_C_bit2(B_config_C[50]),
    .Tile_X0Y2_B_config_C_bit3(B_config_C[51]),
    .Tile_X0Y1_B_config_C_bit0(B_config_C[52]),
    .Tile_X0Y1_B_config_C_bit1(B_config_C[53]),
    .Tile_X0Y1_B_config_C_bit2(B_config_C[54]),
    .Tile_X0Y1_B_config_C_bit3(B_config_C[55]),
    .Tile_X9Y14_Config_accessC_bit0(Config_accessC[0]),
    .Tile_X9Y14_Config_accessC_bit1(Config_accessC[1]),
    .Tile_X9Y14_Config_accessC_bit2(Config_accessC[2]),
    .Tile_X9Y14_Config_accessC_bit3(Config_accessC[3]),
    .Tile_X9Y13_Config_accessC_bit0(Config_accessC[4]),
    .Tile_X9Y13_Config_accessC_bit1(Config_accessC[5]),
    .Tile_X9Y13_Config_accessC_bit2(Config_accessC[6]),
    .Tile_X9Y13_Config_accessC_bit3(Config_accessC[7]),
    .Tile_X9Y12_Config_accessC_bit0(Config_accessC[8]),
    .Tile_X9Y12_Config_accessC_bit1(Config_accessC[9]),
    .Tile_X9Y12_Config_accessC_bit2(Config_accessC[10]),
    .Tile_X9Y12_Config_accessC_bit3(Config_accessC[11]),
    .Tile_X9Y11_Config_accessC_bit0(Config_accessC[12]),
    .Tile_X9Y11_Config_accessC_bit1(Config_accessC[13]),
    .Tile_X9Y11_Config_accessC_bit2(Config_accessC[14]),
    .Tile_X9Y11_Config_accessC_bit3(Config_accessC[15]),
    .Tile_X9Y10_Config_accessC_bit0(Config_accessC[16]),
    .Tile_X9Y10_Config_accessC_bit1(Config_accessC[17]),
    .Tile_X9Y10_Config_accessC_bit2(Config_accessC[18]),
    .Tile_X9Y10_Config_accessC_bit3(Config_accessC[19]),
    .Tile_X9Y9_Config_accessC_bit0(Config_accessC[20]),
    .Tile_X9Y9_Config_accessC_bit1(Config_accessC[21]),
    .Tile_X9Y9_Config_accessC_bit2(Config_accessC[22]),
    .Tile_X9Y9_Config_accessC_bit3(Config_accessC[23]),
    .Tile_X9Y8_Config_accessC_bit0(Config_accessC[24]),
    .Tile_X9Y8_Config_accessC_bit1(Config_accessC[25]),
    .Tile_X9Y8_Config_accessC_bit2(Config_accessC[26]),
    .Tile_X9Y8_Config_accessC_bit3(Config_accessC[27]),
    .Tile_X9Y7_Config_accessC_bit0(Config_accessC[28]),
    .Tile_X9Y7_Config_accessC_bit1(Config_accessC[29]),
    .Tile_X9Y7_Config_accessC_bit2(Config_accessC[30]),
    .Tile_X9Y7_Config_accessC_bit3(Config_accessC[31]),
    .Tile_X9Y6_Config_accessC_bit0(Config_accessC[32]),
    .Tile_X9Y6_Config_accessC_bit1(Config_accessC[33]),
    .Tile_X9Y6_Config_accessC_bit2(Config_accessC[34]),
    .Tile_X9Y6_Config_accessC_bit3(Config_accessC[35]),
    .Tile_X9Y5_Config_accessC_bit0(Config_accessC[36]),
    .Tile_X9Y5_Config_accessC_bit1(Config_accessC[37]),
    .Tile_X9Y5_Config_accessC_bit2(Config_accessC[38]),
    .Tile_X9Y5_Config_accessC_bit3(Config_accessC[39]),
    .Tile_X9Y4_Config_accessC_bit0(Config_accessC[40]),
    .Tile_X9Y4_Config_accessC_bit1(Config_accessC[41]),
    .Tile_X9Y4_Config_accessC_bit2(Config_accessC[42]),
    .Tile_X9Y4_Config_accessC_bit3(Config_accessC[43]),
    .Tile_X9Y3_Config_accessC_bit0(Config_accessC[44]),
    .Tile_X9Y3_Config_accessC_bit1(Config_accessC[45]),
    .Tile_X9Y3_Config_accessC_bit2(Config_accessC[46]),
    .Tile_X9Y3_Config_accessC_bit3(Config_accessC[47]),
    .Tile_X9Y2_Config_accessC_bit0(Config_accessC[48]),
    .Tile_X9Y2_Config_accessC_bit1(Config_accessC[49]),
    .Tile_X9Y2_Config_accessC_bit2(Config_accessC[50]),
    .Tile_X9Y2_Config_accessC_bit3(Config_accessC[51]),
    .Tile_X9Y1_Config_accessC_bit0(Config_accessC[52]),
    .Tile_X9Y1_Config_accessC_bit1(Config_accessC[53]),
    .Tile_X9Y1_Config_accessC_bit2(Config_accessC[54]),
    .Tile_X9Y1_Config_accessC_bit3(Config_accessC[55]),
    .Tile_X9Y14_FAB2RAM_A0_O0(FAB2RAM_A_O[0]),
    .Tile_X9Y14_FAB2RAM_A0_O1(FAB2RAM_A_O[1]),
    .Tile_X9Y14_FAB2RAM_A0_O2(FAB2RAM_A_O[2]),
    .Tile_X9Y14_FAB2RAM_A0_O3(FAB2RAM_A_O[3]),
    .Tile_X9Y14_FAB2RAM_A1_O0(FAB2RAM_A_O[4]),
    .Tile_X9Y14_FAB2RAM_A1_O1(FAB2RAM_A_O[5]),
    .Tile_X9Y14_FAB2RAM_A1_O2(FAB2RAM_A_O[6]),
    .Tile_X9Y14_FAB2RAM_A1_O3(FAB2RAM_A_O[7]),
    .Tile_X9Y13_FAB2RAM_A0_O0(FAB2RAM_A_O[8]),
    .Tile_X9Y13_FAB2RAM_A0_O1(FAB2RAM_A_O[9]),
    .Tile_X9Y13_FAB2RAM_A0_O2(FAB2RAM_A_O[10]),
    .Tile_X9Y13_FAB2RAM_A0_O3(FAB2RAM_A_O[11]),
    .Tile_X9Y13_FAB2RAM_A1_O0(FAB2RAM_A_O[12]),
    .Tile_X9Y13_FAB2RAM_A1_O1(FAB2RAM_A_O[13]),
    .Tile_X9Y13_FAB2RAM_A1_O2(FAB2RAM_A_O[14]),
    .Tile_X9Y13_FAB2RAM_A1_O3(FAB2RAM_A_O[15]),
    .Tile_X9Y12_FAB2RAM_A0_O0(FAB2RAM_A_O[16]),
    .Tile_X9Y12_FAB2RAM_A0_O1(FAB2RAM_A_O[17]),
    .Tile_X9Y12_FAB2RAM_A0_O2(FAB2RAM_A_O[18]),
    .Tile_X9Y12_FAB2RAM_A0_O3(FAB2RAM_A_O[19]),
    .Tile_X9Y12_FAB2RAM_A1_O0(FAB2RAM_A_O[20]),
    .Tile_X9Y12_FAB2RAM_A1_O1(FAB2RAM_A_O[21]),
    .Tile_X9Y12_FAB2RAM_A1_O2(FAB2RAM_A_O[22]),
    .Tile_X9Y12_FAB2RAM_A1_O3(FAB2RAM_A_O[23]),
    .Tile_X9Y11_FAB2RAM_A0_O0(FAB2RAM_A_O[24]),
    .Tile_X9Y11_FAB2RAM_A0_O1(FAB2RAM_A_O[25]),
    .Tile_X9Y11_FAB2RAM_A0_O2(FAB2RAM_A_O[26]),
    .Tile_X9Y11_FAB2RAM_A0_O3(FAB2RAM_A_O[27]),
    .Tile_X9Y11_FAB2RAM_A1_O0(FAB2RAM_A_O[28]),
    .Tile_X9Y11_FAB2RAM_A1_O1(FAB2RAM_A_O[29]),
    .Tile_X9Y11_FAB2RAM_A1_O2(FAB2RAM_A_O[30]),
    .Tile_X9Y11_FAB2RAM_A1_O3(FAB2RAM_A_O[31]),
    .Tile_X9Y10_FAB2RAM_A0_O0(FAB2RAM_A_O[32]),
    .Tile_X9Y10_FAB2RAM_A0_O1(FAB2RAM_A_O[33]),
    .Tile_X9Y10_FAB2RAM_A0_O2(FAB2RAM_A_O[34]),
    .Tile_X9Y10_FAB2RAM_A0_O3(FAB2RAM_A_O[35]),
    .Tile_X9Y10_FAB2RAM_A1_O0(FAB2RAM_A_O[36]),
    .Tile_X9Y10_FAB2RAM_A1_O1(FAB2RAM_A_O[37]),
    .Tile_X9Y10_FAB2RAM_A1_O2(FAB2RAM_A_O[38]),
    .Tile_X9Y10_FAB2RAM_A1_O3(FAB2RAM_A_O[39]),
    .Tile_X9Y9_FAB2RAM_A0_O0(FAB2RAM_A_O[40]),
    .Tile_X9Y9_FAB2RAM_A0_O1(FAB2RAM_A_O[41]),
    .Tile_X9Y9_FAB2RAM_A0_O2(FAB2RAM_A_O[42]),
    .Tile_X9Y9_FAB2RAM_A0_O3(FAB2RAM_A_O[43]),
    .Tile_X9Y9_FAB2RAM_A1_O0(FAB2RAM_A_O[44]),
    .Tile_X9Y9_FAB2RAM_A1_O1(FAB2RAM_A_O[45]),
    .Tile_X9Y9_FAB2RAM_A1_O2(FAB2RAM_A_O[46]),
    .Tile_X9Y9_FAB2RAM_A1_O3(FAB2RAM_A_O[47]),
    .Tile_X9Y8_FAB2RAM_A0_O0(FAB2RAM_A_O[48]),
    .Tile_X9Y8_FAB2RAM_A0_O1(FAB2RAM_A_O[49]),
    .Tile_X9Y8_FAB2RAM_A0_O2(FAB2RAM_A_O[50]),
    .Tile_X9Y8_FAB2RAM_A0_O3(FAB2RAM_A_O[51]),
    .Tile_X9Y8_FAB2RAM_A1_O0(FAB2RAM_A_O[52]),
    .Tile_X9Y8_FAB2RAM_A1_O1(FAB2RAM_A_O[53]),
    .Tile_X9Y8_FAB2RAM_A1_O2(FAB2RAM_A_O[54]),
    .Tile_X9Y8_FAB2RAM_A1_O3(FAB2RAM_A_O[55]),
    .Tile_X9Y7_FAB2RAM_A0_O0(FAB2RAM_A_O[56]),
    .Tile_X9Y7_FAB2RAM_A0_O1(FAB2RAM_A_O[57]),
    .Tile_X9Y7_FAB2RAM_A0_O2(FAB2RAM_A_O[58]),
    .Tile_X9Y7_FAB2RAM_A0_O3(FAB2RAM_A_O[59]),
    .Tile_X9Y7_FAB2RAM_A1_O0(FAB2RAM_A_O[60]),
    .Tile_X9Y7_FAB2RAM_A1_O1(FAB2RAM_A_O[61]),
    .Tile_X9Y7_FAB2RAM_A1_O2(FAB2RAM_A_O[62]),
    .Tile_X9Y7_FAB2RAM_A1_O3(FAB2RAM_A_O[63]),
    .Tile_X9Y6_FAB2RAM_A0_O0(FAB2RAM_A_O[64]),
    .Tile_X9Y6_FAB2RAM_A0_O1(FAB2RAM_A_O[65]),
    .Tile_X9Y6_FAB2RAM_A0_O2(FAB2RAM_A_O[66]),
    .Tile_X9Y6_FAB2RAM_A0_O3(FAB2RAM_A_O[67]),
    .Tile_X9Y6_FAB2RAM_A1_O0(FAB2RAM_A_O[68]),
    .Tile_X9Y6_FAB2RAM_A1_O1(FAB2RAM_A_O[69]),
    .Tile_X9Y6_FAB2RAM_A1_O2(FAB2RAM_A_O[70]),
    .Tile_X9Y6_FAB2RAM_A1_O3(FAB2RAM_A_O[71]),
    .Tile_X9Y5_FAB2RAM_A0_O0(FAB2RAM_A_O[72]),
    .Tile_X9Y5_FAB2RAM_A0_O1(FAB2RAM_A_O[73]),
    .Tile_X9Y5_FAB2RAM_A0_O2(FAB2RAM_A_O[74]),
    .Tile_X9Y5_FAB2RAM_A0_O3(FAB2RAM_A_O[75]),
    .Tile_X9Y5_FAB2RAM_A1_O0(FAB2RAM_A_O[76]),
    .Tile_X9Y5_FAB2RAM_A1_O1(FAB2RAM_A_O[77]),
    .Tile_X9Y5_FAB2RAM_A1_O2(FAB2RAM_A_O[78]),
    .Tile_X9Y5_FAB2RAM_A1_O3(FAB2RAM_A_O[79]),
    .Tile_X9Y4_FAB2RAM_A0_O0(FAB2RAM_A_O[80]),
    .Tile_X9Y4_FAB2RAM_A0_O1(FAB2RAM_A_O[81]),
    .Tile_X9Y4_FAB2RAM_A0_O2(FAB2RAM_A_O[82]),
    .Tile_X9Y4_FAB2RAM_A0_O3(FAB2RAM_A_O[83]),
    .Tile_X9Y4_FAB2RAM_A1_O0(FAB2RAM_A_O[84]),
    .Tile_X9Y4_FAB2RAM_A1_O1(FAB2RAM_A_O[85]),
    .Tile_X9Y4_FAB2RAM_A1_O2(FAB2RAM_A_O[86]),
    .Tile_X9Y4_FAB2RAM_A1_O3(FAB2RAM_A_O[87]),
    .Tile_X9Y3_FAB2RAM_A0_O0(FAB2RAM_A_O[88]),
    .Tile_X9Y3_FAB2RAM_A0_O1(FAB2RAM_A_O[89]),
    .Tile_X9Y3_FAB2RAM_A0_O2(FAB2RAM_A_O[90]),
    .Tile_X9Y3_FAB2RAM_A0_O3(FAB2RAM_A_O[91]),
    .Tile_X9Y3_FAB2RAM_A1_O0(FAB2RAM_A_O[92]),
    .Tile_X9Y3_FAB2RAM_A1_O1(FAB2RAM_A_O[93]),
    .Tile_X9Y3_FAB2RAM_A1_O2(FAB2RAM_A_O[94]),
    .Tile_X9Y3_FAB2RAM_A1_O3(FAB2RAM_A_O[95]),
    .Tile_X9Y2_FAB2RAM_A0_O0(FAB2RAM_A_O[96]),
    .Tile_X9Y2_FAB2RAM_A0_O1(FAB2RAM_A_O[97]),
    .Tile_X9Y2_FAB2RAM_A0_O2(FAB2RAM_A_O[98]),
    .Tile_X9Y2_FAB2RAM_A0_O3(FAB2RAM_A_O[99]),
    .Tile_X9Y2_FAB2RAM_A1_O0(FAB2RAM_A_O[100]),
    .Tile_X9Y2_FAB2RAM_A1_O1(FAB2RAM_A_O[101]),
    .Tile_X9Y2_FAB2RAM_A1_O2(FAB2RAM_A_O[102]),
    .Tile_X9Y2_FAB2RAM_A1_O3(FAB2RAM_A_O[103]),
    .Tile_X9Y1_FAB2RAM_A0_O0(FAB2RAM_A_O[104]),
    .Tile_X9Y1_FAB2RAM_A0_O1(FAB2RAM_A_O[105]),
    .Tile_X9Y1_FAB2RAM_A0_O2(FAB2RAM_A_O[106]),
    .Tile_X9Y1_FAB2RAM_A0_O3(FAB2RAM_A_O[107]),
    .Tile_X9Y1_FAB2RAM_A1_O0(FAB2RAM_A_O[108]),
    .Tile_X9Y1_FAB2RAM_A1_O1(FAB2RAM_A_O[109]),
    .Tile_X9Y1_FAB2RAM_A1_O2(FAB2RAM_A_O[110]),
    .Tile_X9Y1_FAB2RAM_A1_O3(FAB2RAM_A_O[111]),
    .Tile_X9Y14_FAB2RAM_C_O0(FAB2RAM_C_O[0]),
    .Tile_X9Y14_FAB2RAM_C_O1(FAB2RAM_C_O[1]),
    .Tile_X9Y14_FAB2RAM_C_O2(FAB2RAM_C_O[2]),
    .Tile_X9Y14_FAB2RAM_C_O3(FAB2RAM_C_O[3]),
    .Tile_X9Y13_FAB2RAM_C_O0(FAB2RAM_C_O[4]),
    .Tile_X9Y13_FAB2RAM_C_O1(FAB2RAM_C_O[5]),
    .Tile_X9Y13_FAB2RAM_C_O2(FAB2RAM_C_O[6]),
    .Tile_X9Y13_FAB2RAM_C_O3(FAB2RAM_C_O[7]),
    .Tile_X9Y12_FAB2RAM_C_O0(FAB2RAM_C_O[8]),
    .Tile_X9Y12_FAB2RAM_C_O1(FAB2RAM_C_O[9]),
    .Tile_X9Y12_FAB2RAM_C_O2(FAB2RAM_C_O[10]),
    .Tile_X9Y12_FAB2RAM_C_O3(FAB2RAM_C_O[11]),
    .Tile_X9Y11_FAB2RAM_C_O0(FAB2RAM_C_O[12]),
    .Tile_X9Y11_FAB2RAM_C_O1(FAB2RAM_C_O[13]),
    .Tile_X9Y11_FAB2RAM_C_O2(FAB2RAM_C_O[14]),
    .Tile_X9Y11_FAB2RAM_C_O3(FAB2RAM_C_O[15]),
    .Tile_X9Y10_FAB2RAM_C_O0(FAB2RAM_C_O[16]),
    .Tile_X9Y10_FAB2RAM_C_O1(FAB2RAM_C_O[17]),
    .Tile_X9Y10_FAB2RAM_C_O2(FAB2RAM_C_O[18]),
    .Tile_X9Y10_FAB2RAM_C_O3(FAB2RAM_C_O[19]),
    .Tile_X9Y9_FAB2RAM_C_O0(FAB2RAM_C_O[20]),
    .Tile_X9Y9_FAB2RAM_C_O1(FAB2RAM_C_O[21]),
    .Tile_X9Y9_FAB2RAM_C_O2(FAB2RAM_C_O[22]),
    .Tile_X9Y9_FAB2RAM_C_O3(FAB2RAM_C_O[23]),
    .Tile_X9Y8_FAB2RAM_C_O0(FAB2RAM_C_O[24]),
    .Tile_X9Y8_FAB2RAM_C_O1(FAB2RAM_C_O[25]),
    .Tile_X9Y8_FAB2RAM_C_O2(FAB2RAM_C_O[26]),
    .Tile_X9Y8_FAB2RAM_C_O3(FAB2RAM_C_O[27]),
    .Tile_X9Y7_FAB2RAM_C_O0(FAB2RAM_C_O[28]),
    .Tile_X9Y7_FAB2RAM_C_O1(FAB2RAM_C_O[29]),
    .Tile_X9Y7_FAB2RAM_C_O2(FAB2RAM_C_O[30]),
    .Tile_X9Y7_FAB2RAM_C_O3(FAB2RAM_C_O[31]),
    .Tile_X9Y6_FAB2RAM_C_O0(FAB2RAM_C_O[32]),
    .Tile_X9Y6_FAB2RAM_C_O1(FAB2RAM_C_O[33]),
    .Tile_X9Y6_FAB2RAM_C_O2(FAB2RAM_C_O[34]),
    .Tile_X9Y6_FAB2RAM_C_O3(FAB2RAM_C_O[35]),
    .Tile_X9Y5_FAB2RAM_C_O0(FAB2RAM_C_O[36]),
    .Tile_X9Y5_FAB2RAM_C_O1(FAB2RAM_C_O[37]),
    .Tile_X9Y5_FAB2RAM_C_O2(FAB2RAM_C_O[38]),
    .Tile_X9Y5_FAB2RAM_C_O3(FAB2RAM_C_O[39]),
    .Tile_X9Y4_FAB2RAM_C_O0(FAB2RAM_C_O[40]),
    .Tile_X9Y4_FAB2RAM_C_O1(FAB2RAM_C_O[41]),
    .Tile_X9Y4_FAB2RAM_C_O2(FAB2RAM_C_O[42]),
    .Tile_X9Y4_FAB2RAM_C_O3(FAB2RAM_C_O[43]),
    .Tile_X9Y3_FAB2RAM_C_O0(FAB2RAM_C_O[44]),
    .Tile_X9Y3_FAB2RAM_C_O1(FAB2RAM_C_O[45]),
    .Tile_X9Y3_FAB2RAM_C_O2(FAB2RAM_C_O[46]),
    .Tile_X9Y3_FAB2RAM_C_O3(FAB2RAM_C_O[47]),
    .Tile_X9Y2_FAB2RAM_C_O0(FAB2RAM_C_O[48]),
    .Tile_X9Y2_FAB2RAM_C_O1(FAB2RAM_C_O[49]),
    .Tile_X9Y2_FAB2RAM_C_O2(FAB2RAM_C_O[50]),
    .Tile_X9Y2_FAB2RAM_C_O3(FAB2RAM_C_O[51]),
    .Tile_X9Y1_FAB2RAM_C_O0(FAB2RAM_C_O[52]),
    .Tile_X9Y1_FAB2RAM_C_O1(FAB2RAM_C_O[53]),
    .Tile_X9Y1_FAB2RAM_C_O2(FAB2RAM_C_O[54]),
    .Tile_X9Y1_FAB2RAM_C_O3(FAB2RAM_C_O[55]),
    .Tile_X9Y14_FAB2RAM_D0_O0(FAB2RAM_D_O[0]),
    .Tile_X9Y14_FAB2RAM_D0_O1(FAB2RAM_D_O[1]),
    .Tile_X9Y14_FAB2RAM_D0_O2(FAB2RAM_D_O[2]),
    .Tile_X9Y14_FAB2RAM_D0_O3(FAB2RAM_D_O[3]),
    .Tile_X9Y14_FAB2RAM_D1_O0(FAB2RAM_D_O[4]),
    .Tile_X9Y14_FAB2RAM_D1_O1(FAB2RAM_D_O[5]),
    .Tile_X9Y14_FAB2RAM_D1_O2(FAB2RAM_D_O[6]),
    .Tile_X9Y14_FAB2RAM_D1_O3(FAB2RAM_D_O[7]),
    .Tile_X9Y14_FAB2RAM_D2_O0(FAB2RAM_D_O[8]),
    .Tile_X9Y14_FAB2RAM_D2_O1(FAB2RAM_D_O[9]),
    .Tile_X9Y14_FAB2RAM_D2_O2(FAB2RAM_D_O[10]),
    .Tile_X9Y14_FAB2RAM_D2_O3(FAB2RAM_D_O[11]),
    .Tile_X9Y14_FAB2RAM_D3_O0(FAB2RAM_D_O[12]),
    .Tile_X9Y14_FAB2RAM_D3_O1(FAB2RAM_D_O[13]),
    .Tile_X9Y14_FAB2RAM_D3_O2(FAB2RAM_D_O[14]),
    .Tile_X9Y14_FAB2RAM_D3_O3(FAB2RAM_D_O[15]),
    .Tile_X9Y13_FAB2RAM_D0_O0(FAB2RAM_D_O[16]),
    .Tile_X9Y13_FAB2RAM_D0_O1(FAB2RAM_D_O[17]),
    .Tile_X9Y13_FAB2RAM_D0_O2(FAB2RAM_D_O[18]),
    .Tile_X9Y13_FAB2RAM_D0_O3(FAB2RAM_D_O[19]),
    .Tile_X9Y13_FAB2RAM_D1_O0(FAB2RAM_D_O[20]),
    .Tile_X9Y13_FAB2RAM_D1_O1(FAB2RAM_D_O[21]),
    .Tile_X9Y13_FAB2RAM_D1_O2(FAB2RAM_D_O[22]),
    .Tile_X9Y13_FAB2RAM_D1_O3(FAB2RAM_D_O[23]),
    .Tile_X9Y13_FAB2RAM_D2_O0(FAB2RAM_D_O[24]),
    .Tile_X9Y13_FAB2RAM_D2_O1(FAB2RAM_D_O[25]),
    .Tile_X9Y13_FAB2RAM_D2_O2(FAB2RAM_D_O[26]),
    .Tile_X9Y13_FAB2RAM_D2_O3(FAB2RAM_D_O[27]),
    .Tile_X9Y13_FAB2RAM_D3_O0(FAB2RAM_D_O[28]),
    .Tile_X9Y13_FAB2RAM_D3_O1(FAB2RAM_D_O[29]),
    .Tile_X9Y13_FAB2RAM_D3_O2(FAB2RAM_D_O[30]),
    .Tile_X9Y13_FAB2RAM_D3_O3(FAB2RAM_D_O[31]),
    .Tile_X9Y12_FAB2RAM_D0_O0(FAB2RAM_D_O[32]),
    .Tile_X9Y12_FAB2RAM_D0_O1(FAB2RAM_D_O[33]),
    .Tile_X9Y12_FAB2RAM_D0_O2(FAB2RAM_D_O[34]),
    .Tile_X9Y12_FAB2RAM_D0_O3(FAB2RAM_D_O[35]),
    .Tile_X9Y12_FAB2RAM_D1_O0(FAB2RAM_D_O[36]),
    .Tile_X9Y12_FAB2RAM_D1_O1(FAB2RAM_D_O[37]),
    .Tile_X9Y12_FAB2RAM_D1_O2(FAB2RAM_D_O[38]),
    .Tile_X9Y12_FAB2RAM_D1_O3(FAB2RAM_D_O[39]),
    .Tile_X9Y12_FAB2RAM_D2_O0(FAB2RAM_D_O[40]),
    .Tile_X9Y12_FAB2RAM_D2_O1(FAB2RAM_D_O[41]),
    .Tile_X9Y12_FAB2RAM_D2_O2(FAB2RAM_D_O[42]),
    .Tile_X9Y12_FAB2RAM_D2_O3(FAB2RAM_D_O[43]),
    .Tile_X9Y12_FAB2RAM_D3_O0(FAB2RAM_D_O[44]),
    .Tile_X9Y12_FAB2RAM_D3_O1(FAB2RAM_D_O[45]),
    .Tile_X9Y12_FAB2RAM_D3_O2(FAB2RAM_D_O[46]),
    .Tile_X9Y12_FAB2RAM_D3_O3(FAB2RAM_D_O[47]),
    .Tile_X9Y11_FAB2RAM_D0_O0(FAB2RAM_D_O[48]),
    .Tile_X9Y11_FAB2RAM_D0_O1(FAB2RAM_D_O[49]),
    .Tile_X9Y11_FAB2RAM_D0_O2(FAB2RAM_D_O[50]),
    .Tile_X9Y11_FAB2RAM_D0_O3(FAB2RAM_D_O[51]),
    .Tile_X9Y11_FAB2RAM_D1_O0(FAB2RAM_D_O[52]),
    .Tile_X9Y11_FAB2RAM_D1_O1(FAB2RAM_D_O[53]),
    .Tile_X9Y11_FAB2RAM_D1_O2(FAB2RAM_D_O[54]),
    .Tile_X9Y11_FAB2RAM_D1_O3(FAB2RAM_D_O[55]),
    .Tile_X9Y11_FAB2RAM_D2_O0(FAB2RAM_D_O[56]),
    .Tile_X9Y11_FAB2RAM_D2_O1(FAB2RAM_D_O[57]),
    .Tile_X9Y11_FAB2RAM_D2_O2(FAB2RAM_D_O[58]),
    .Tile_X9Y11_FAB2RAM_D2_O3(FAB2RAM_D_O[59]),
    .Tile_X9Y11_FAB2RAM_D3_O0(FAB2RAM_D_O[60]),
    .Tile_X9Y11_FAB2RAM_D3_O1(FAB2RAM_D_O[61]),
    .Tile_X9Y11_FAB2RAM_D3_O2(FAB2RAM_D_O[62]),
    .Tile_X9Y11_FAB2RAM_D3_O3(FAB2RAM_D_O[63]),
    .Tile_X9Y10_FAB2RAM_D0_O0(FAB2RAM_D_O[64]),
    .Tile_X9Y10_FAB2RAM_D0_O1(FAB2RAM_D_O[65]),
    .Tile_X9Y10_FAB2RAM_D0_O2(FAB2RAM_D_O[66]),
    .Tile_X9Y10_FAB2RAM_D0_O3(FAB2RAM_D_O[67]),
    .Tile_X9Y10_FAB2RAM_D1_O0(FAB2RAM_D_O[68]),
    .Tile_X9Y10_FAB2RAM_D1_O1(FAB2RAM_D_O[69]),
    .Tile_X9Y10_FAB2RAM_D1_O2(FAB2RAM_D_O[70]),
    .Tile_X9Y10_FAB2RAM_D1_O3(FAB2RAM_D_O[71]),
    .Tile_X9Y10_FAB2RAM_D2_O0(FAB2RAM_D_O[72]),
    .Tile_X9Y10_FAB2RAM_D2_O1(FAB2RAM_D_O[73]),
    .Tile_X9Y10_FAB2RAM_D2_O2(FAB2RAM_D_O[74]),
    .Tile_X9Y10_FAB2RAM_D2_O3(FAB2RAM_D_O[75]),
    .Tile_X9Y10_FAB2RAM_D3_O0(FAB2RAM_D_O[76]),
    .Tile_X9Y10_FAB2RAM_D3_O1(FAB2RAM_D_O[77]),
    .Tile_X9Y10_FAB2RAM_D3_O2(FAB2RAM_D_O[78]),
    .Tile_X9Y10_FAB2RAM_D3_O3(FAB2RAM_D_O[79]),
    .Tile_X9Y9_FAB2RAM_D0_O0(FAB2RAM_D_O[80]),
    .Tile_X9Y9_FAB2RAM_D0_O1(FAB2RAM_D_O[81]),
    .Tile_X9Y9_FAB2RAM_D0_O2(FAB2RAM_D_O[82]),
    .Tile_X9Y9_FAB2RAM_D0_O3(FAB2RAM_D_O[83]),
    .Tile_X9Y9_FAB2RAM_D1_O0(FAB2RAM_D_O[84]),
    .Tile_X9Y9_FAB2RAM_D1_O1(FAB2RAM_D_O[85]),
    .Tile_X9Y9_FAB2RAM_D1_O2(FAB2RAM_D_O[86]),
    .Tile_X9Y9_FAB2RAM_D1_O3(FAB2RAM_D_O[87]),
    .Tile_X9Y9_FAB2RAM_D2_O0(FAB2RAM_D_O[88]),
    .Tile_X9Y9_FAB2RAM_D2_O1(FAB2RAM_D_O[89]),
    .Tile_X9Y9_FAB2RAM_D2_O2(FAB2RAM_D_O[90]),
    .Tile_X9Y9_FAB2RAM_D2_O3(FAB2RAM_D_O[91]),
    .Tile_X9Y9_FAB2RAM_D3_O0(FAB2RAM_D_O[92]),
    .Tile_X9Y9_FAB2RAM_D3_O1(FAB2RAM_D_O[93]),
    .Tile_X9Y9_FAB2RAM_D3_O2(FAB2RAM_D_O[94]),
    .Tile_X9Y9_FAB2RAM_D3_O3(FAB2RAM_D_O[95]),
    .Tile_X9Y8_FAB2RAM_D0_O0(FAB2RAM_D_O[96]),
    .Tile_X9Y8_FAB2RAM_D0_O1(FAB2RAM_D_O[97]),
    .Tile_X9Y8_FAB2RAM_D0_O2(FAB2RAM_D_O[98]),
    .Tile_X9Y8_FAB2RAM_D0_O3(FAB2RAM_D_O[99]),
    .Tile_X9Y8_FAB2RAM_D1_O0(FAB2RAM_D_O[100]),
    .Tile_X9Y8_FAB2RAM_D1_O1(FAB2RAM_D_O[101]),
    .Tile_X9Y8_FAB2RAM_D1_O2(FAB2RAM_D_O[102]),
    .Tile_X9Y8_FAB2RAM_D1_O3(FAB2RAM_D_O[103]),
    .Tile_X9Y8_FAB2RAM_D2_O0(FAB2RAM_D_O[104]),
    .Tile_X9Y8_FAB2RAM_D2_O1(FAB2RAM_D_O[105]),
    .Tile_X9Y8_FAB2RAM_D2_O2(FAB2RAM_D_O[106]),
    .Tile_X9Y8_FAB2RAM_D2_O3(FAB2RAM_D_O[107]),
    .Tile_X9Y8_FAB2RAM_D3_O0(FAB2RAM_D_O[108]),
    .Tile_X9Y8_FAB2RAM_D3_O1(FAB2RAM_D_O[109]),
    .Tile_X9Y8_FAB2RAM_D3_O2(FAB2RAM_D_O[110]),
    .Tile_X9Y8_FAB2RAM_D3_O3(FAB2RAM_D_O[111]),
    .Tile_X9Y7_FAB2RAM_D0_O0(FAB2RAM_D_O[112]),
    .Tile_X9Y7_FAB2RAM_D0_O1(FAB2RAM_D_O[113]),
    .Tile_X9Y7_FAB2RAM_D0_O2(FAB2RAM_D_O[114]),
    .Tile_X9Y7_FAB2RAM_D0_O3(FAB2RAM_D_O[115]),
    .Tile_X9Y7_FAB2RAM_D1_O0(FAB2RAM_D_O[116]),
    .Tile_X9Y7_FAB2RAM_D1_O1(FAB2RAM_D_O[117]),
    .Tile_X9Y7_FAB2RAM_D1_O2(FAB2RAM_D_O[118]),
    .Tile_X9Y7_FAB2RAM_D1_O3(FAB2RAM_D_O[119]),
    .Tile_X9Y7_FAB2RAM_D2_O0(FAB2RAM_D_O[120]),
    .Tile_X9Y7_FAB2RAM_D2_O1(FAB2RAM_D_O[121]),
    .Tile_X9Y7_FAB2RAM_D2_O2(FAB2RAM_D_O[122]),
    .Tile_X9Y7_FAB2RAM_D2_O3(FAB2RAM_D_O[123]),
    .Tile_X9Y7_FAB2RAM_D3_O0(FAB2RAM_D_O[124]),
    .Tile_X9Y7_FAB2RAM_D3_O1(FAB2RAM_D_O[125]),
    .Tile_X9Y7_FAB2RAM_D3_O2(FAB2RAM_D_O[126]),
    .Tile_X9Y7_FAB2RAM_D3_O3(FAB2RAM_D_O[127]),
    .Tile_X9Y6_FAB2RAM_D0_O0(FAB2RAM_D_O[128]),
    .Tile_X9Y6_FAB2RAM_D0_O1(FAB2RAM_D_O[129]),
    .Tile_X9Y6_FAB2RAM_D0_O2(FAB2RAM_D_O[130]),
    .Tile_X9Y6_FAB2RAM_D0_O3(FAB2RAM_D_O[131]),
    .Tile_X9Y6_FAB2RAM_D1_O0(FAB2RAM_D_O[132]),
    .Tile_X9Y6_FAB2RAM_D1_O1(FAB2RAM_D_O[133]),
    .Tile_X9Y6_FAB2RAM_D1_O2(FAB2RAM_D_O[134]),
    .Tile_X9Y6_FAB2RAM_D1_O3(FAB2RAM_D_O[135]),
    .Tile_X9Y6_FAB2RAM_D2_O0(FAB2RAM_D_O[136]),
    .Tile_X9Y6_FAB2RAM_D2_O1(FAB2RAM_D_O[137]),
    .Tile_X9Y6_FAB2RAM_D2_O2(FAB2RAM_D_O[138]),
    .Tile_X9Y6_FAB2RAM_D2_O3(FAB2RAM_D_O[139]),
    .Tile_X9Y6_FAB2RAM_D3_O0(FAB2RAM_D_O[140]),
    .Tile_X9Y6_FAB2RAM_D3_O1(FAB2RAM_D_O[141]),
    .Tile_X9Y6_FAB2RAM_D3_O2(FAB2RAM_D_O[142]),
    .Tile_X9Y6_FAB2RAM_D3_O3(FAB2RAM_D_O[143]),
    .Tile_X9Y5_FAB2RAM_D0_O0(FAB2RAM_D_O[144]),
    .Tile_X9Y5_FAB2RAM_D0_O1(FAB2RAM_D_O[145]),
    .Tile_X9Y5_FAB2RAM_D0_O2(FAB2RAM_D_O[146]),
    .Tile_X9Y5_FAB2RAM_D0_O3(FAB2RAM_D_O[147]),
    .Tile_X9Y5_FAB2RAM_D1_O0(FAB2RAM_D_O[148]),
    .Tile_X9Y5_FAB2RAM_D1_O1(FAB2RAM_D_O[149]),
    .Tile_X9Y5_FAB2RAM_D1_O2(FAB2RAM_D_O[150]),
    .Tile_X9Y5_FAB2RAM_D1_O3(FAB2RAM_D_O[151]),
    .Tile_X9Y5_FAB2RAM_D2_O0(FAB2RAM_D_O[152]),
    .Tile_X9Y5_FAB2RAM_D2_O1(FAB2RAM_D_O[153]),
    .Tile_X9Y5_FAB2RAM_D2_O2(FAB2RAM_D_O[154]),
    .Tile_X9Y5_FAB2RAM_D2_O3(FAB2RAM_D_O[155]),
    .Tile_X9Y5_FAB2RAM_D3_O0(FAB2RAM_D_O[156]),
    .Tile_X9Y5_FAB2RAM_D3_O1(FAB2RAM_D_O[157]),
    .Tile_X9Y5_FAB2RAM_D3_O2(FAB2RAM_D_O[158]),
    .Tile_X9Y5_FAB2RAM_D3_O3(FAB2RAM_D_O[159]),
    .Tile_X9Y4_FAB2RAM_D0_O0(FAB2RAM_D_O[160]),
    .Tile_X9Y4_FAB2RAM_D0_O1(FAB2RAM_D_O[161]),
    .Tile_X9Y4_FAB2RAM_D0_O2(FAB2RAM_D_O[162]),
    .Tile_X9Y4_FAB2RAM_D0_O3(FAB2RAM_D_O[163]),
    .Tile_X9Y4_FAB2RAM_D1_O0(FAB2RAM_D_O[164]),
    .Tile_X9Y4_FAB2RAM_D1_O1(FAB2RAM_D_O[165]),
    .Tile_X9Y4_FAB2RAM_D1_O2(FAB2RAM_D_O[166]),
    .Tile_X9Y4_FAB2RAM_D1_O3(FAB2RAM_D_O[167]),
    .Tile_X9Y4_FAB2RAM_D2_O0(FAB2RAM_D_O[168]),
    .Tile_X9Y4_FAB2RAM_D2_O1(FAB2RAM_D_O[169]),
    .Tile_X9Y4_FAB2RAM_D2_O2(FAB2RAM_D_O[170]),
    .Tile_X9Y4_FAB2RAM_D2_O3(FAB2RAM_D_O[171]),
    .Tile_X9Y4_FAB2RAM_D3_O0(FAB2RAM_D_O[172]),
    .Tile_X9Y4_FAB2RAM_D3_O1(FAB2RAM_D_O[173]),
    .Tile_X9Y4_FAB2RAM_D3_O2(FAB2RAM_D_O[174]),
    .Tile_X9Y4_FAB2RAM_D3_O3(FAB2RAM_D_O[175]),
    .Tile_X9Y3_FAB2RAM_D0_O0(FAB2RAM_D_O[176]),
    .Tile_X9Y3_FAB2RAM_D0_O1(FAB2RAM_D_O[177]),
    .Tile_X9Y3_FAB2RAM_D0_O2(FAB2RAM_D_O[178]),
    .Tile_X9Y3_FAB2RAM_D0_O3(FAB2RAM_D_O[179]),
    .Tile_X9Y3_FAB2RAM_D1_O0(FAB2RAM_D_O[180]),
    .Tile_X9Y3_FAB2RAM_D1_O1(FAB2RAM_D_O[181]),
    .Tile_X9Y3_FAB2RAM_D1_O2(FAB2RAM_D_O[182]),
    .Tile_X9Y3_FAB2RAM_D1_O3(FAB2RAM_D_O[183]),
    .Tile_X9Y3_FAB2RAM_D2_O0(FAB2RAM_D_O[184]),
    .Tile_X9Y3_FAB2RAM_D2_O1(FAB2RAM_D_O[185]),
    .Tile_X9Y3_FAB2RAM_D2_O2(FAB2RAM_D_O[186]),
    .Tile_X9Y3_FAB2RAM_D2_O3(FAB2RAM_D_O[187]),
    .Tile_X9Y3_FAB2RAM_D3_O0(FAB2RAM_D_O[188]),
    .Tile_X9Y3_FAB2RAM_D3_O1(FAB2RAM_D_O[189]),
    .Tile_X9Y3_FAB2RAM_D3_O2(FAB2RAM_D_O[190]),
    .Tile_X9Y3_FAB2RAM_D3_O3(FAB2RAM_D_O[191]),
    .Tile_X9Y2_FAB2RAM_D0_O0(FAB2RAM_D_O[192]),
    .Tile_X9Y2_FAB2RAM_D0_O1(FAB2RAM_D_O[193]),
    .Tile_X9Y2_FAB2RAM_D0_O2(FAB2RAM_D_O[194]),
    .Tile_X9Y2_FAB2RAM_D0_O3(FAB2RAM_D_O[195]),
    .Tile_X9Y2_FAB2RAM_D1_O0(FAB2RAM_D_O[196]),
    .Tile_X9Y2_FAB2RAM_D1_O1(FAB2RAM_D_O[197]),
    .Tile_X9Y2_FAB2RAM_D1_O2(FAB2RAM_D_O[198]),
    .Tile_X9Y2_FAB2RAM_D1_O3(FAB2RAM_D_O[199]),
    .Tile_X9Y2_FAB2RAM_D2_O0(FAB2RAM_D_O[200]),
    .Tile_X9Y2_FAB2RAM_D2_O1(FAB2RAM_D_O[201]),
    .Tile_X9Y2_FAB2RAM_D2_O2(FAB2RAM_D_O[202]),
    .Tile_X9Y2_FAB2RAM_D2_O3(FAB2RAM_D_O[203]),
    .Tile_X9Y2_FAB2RAM_D3_O0(FAB2RAM_D_O[204]),
    .Tile_X9Y2_FAB2RAM_D3_O1(FAB2RAM_D_O[205]),
    .Tile_X9Y2_FAB2RAM_D3_O2(FAB2RAM_D_O[206]),
    .Tile_X9Y2_FAB2RAM_D3_O3(FAB2RAM_D_O[207]),
    .Tile_X9Y1_FAB2RAM_D0_O0(FAB2RAM_D_O[208]),
    .Tile_X9Y1_FAB2RAM_D0_O1(FAB2RAM_D_O[209]),
    .Tile_X9Y1_FAB2RAM_D0_O2(FAB2RAM_D_O[210]),
    .Tile_X9Y1_FAB2RAM_D0_O3(FAB2RAM_D_O[211]),
    .Tile_X9Y1_FAB2RAM_D1_O0(FAB2RAM_D_O[212]),
    .Tile_X9Y1_FAB2RAM_D1_O1(FAB2RAM_D_O[213]),
    .Tile_X9Y1_FAB2RAM_D1_O2(FAB2RAM_D_O[214]),
    .Tile_X9Y1_FAB2RAM_D1_O3(FAB2RAM_D_O[215]),
    .Tile_X9Y1_FAB2RAM_D2_O0(FAB2RAM_D_O[216]),
    .Tile_X9Y1_FAB2RAM_D2_O1(FAB2RAM_D_O[217]),
    .Tile_X9Y1_FAB2RAM_D2_O2(FAB2RAM_D_O[218]),
    .Tile_X9Y1_FAB2RAM_D2_O3(FAB2RAM_D_O[219]),
    .Tile_X9Y1_FAB2RAM_D3_O0(FAB2RAM_D_O[220]),
    .Tile_X9Y1_FAB2RAM_D3_O1(FAB2RAM_D_O[221]),
    .Tile_X9Y1_FAB2RAM_D3_O2(FAB2RAM_D_O[222]),
    .Tile_X9Y1_FAB2RAM_D3_O3(FAB2RAM_D_O[223]),
    .Tile_X0Y14_B_I_top(I_top[0]),
    .Tile_X0Y14_A_I_top(I_top[1]),
    .Tile_X0Y13_B_I_top(I_top[2]),
    .Tile_X0Y13_A_I_top(I_top[3]),
    .Tile_X0Y12_B_I_top(I_top[4]),
    .Tile_X0Y12_A_I_top(I_top[5]),
    .Tile_X0Y11_B_I_top(I_top[6]),
    .Tile_X0Y11_A_I_top(I_top[7]),
    .Tile_X0Y10_B_I_top(I_top[8]),
    .Tile_X0Y10_A_I_top(I_top[9]),
    .Tile_X0Y9_B_I_top(I_top[10]),
    .Tile_X0Y9_A_I_top(I_top[11]),
    .Tile_X0Y8_B_I_top(I_top[12]),
    .Tile_X0Y8_A_I_top(I_top[13]),
    .Tile_X0Y7_B_I_top(I_top[14]),
    .Tile_X0Y7_A_I_top(I_top[15]),
    .Tile_X0Y6_B_I_top(I_top[16]),
    .Tile_X0Y6_A_I_top(I_top[17]),
    .Tile_X0Y5_B_I_top(I_top[18]),
    .Tile_X0Y5_A_I_top(I_top[19]),
    .Tile_X0Y4_B_I_top(I_top[20]),
    .Tile_X0Y4_A_I_top(I_top[21]),
    .Tile_X0Y3_B_I_top(I_top[22]),
    .Tile_X0Y3_A_I_top(I_top[23]),
    .Tile_X0Y2_B_I_top(I_top[24]),
    .Tile_X0Y2_A_I_top(I_top[25]),
    .Tile_X0Y1_B_I_top(I_top[26]),
    .Tile_X0Y1_A_I_top(I_top[27]),
    .Tile_X0Y14_B_O_top(O_top[0]),
    .Tile_X0Y14_A_O_top(O_top[1]),
    .Tile_X0Y13_B_O_top(O_top[2]),
    .Tile_X0Y13_A_O_top(O_top[3]),
    .Tile_X0Y12_B_O_top(O_top[4]),
    .Tile_X0Y12_A_O_top(O_top[5]),
    .Tile_X0Y11_B_O_top(O_top[6]),
    .Tile_X0Y11_A_O_top(O_top[7]),
    .Tile_X0Y10_B_O_top(O_top[8]),
    .Tile_X0Y10_A_O_top(O_top[9]),
    .Tile_X0Y9_B_O_top(O_top[10]),
    .Tile_X0Y9_A_O_top(O_top[11]),
    .Tile_X0Y8_B_O_top(O_top[12]),
    .Tile_X0Y8_A_O_top(O_top[13]),
    .Tile_X0Y7_B_O_top(O_top[14]),
    .Tile_X0Y7_A_O_top(O_top[15]),
    .Tile_X0Y6_B_O_top(O_top[16]),
    .Tile_X0Y6_A_O_top(O_top[17]),
    .Tile_X0Y5_B_O_top(O_top[18]),
    .Tile_X0Y5_A_O_top(O_top[19]),
    .Tile_X0Y4_B_O_top(O_top[20]),
    .Tile_X0Y4_A_O_top(O_top[21]),
    .Tile_X0Y3_B_O_top(O_top[22]),
    .Tile_X0Y3_A_O_top(O_top[23]),
    .Tile_X0Y2_B_O_top(O_top[24]),
    .Tile_X0Y2_A_O_top(O_top[25]),
    .Tile_X0Y1_B_O_top(O_top[26]),
    .Tile_X0Y1_A_O_top(O_top[27]),
    .Tile_X9Y14_RAM2FAB_D0_I0(RAM2FAB_D_I[0]),
    .Tile_X9Y14_RAM2FAB_D0_I1(RAM2FAB_D_I[1]),
    .Tile_X9Y14_RAM2FAB_D0_I2(RAM2FAB_D_I[2]),
    .Tile_X9Y14_RAM2FAB_D0_I3(RAM2FAB_D_I[3]),
    .Tile_X9Y14_RAM2FAB_D1_I0(RAM2FAB_D_I[4]),
    .Tile_X9Y14_RAM2FAB_D1_I1(RAM2FAB_D_I[5]),
    .Tile_X9Y14_RAM2FAB_D1_I2(RAM2FAB_D_I[6]),
    .Tile_X9Y14_RAM2FAB_D1_I3(RAM2FAB_D_I[7]),
    .Tile_X9Y14_RAM2FAB_D2_I0(RAM2FAB_D_I[8]),
    .Tile_X9Y14_RAM2FAB_D2_I1(RAM2FAB_D_I[9]),
    .Tile_X9Y14_RAM2FAB_D2_I2(RAM2FAB_D_I[10]),
    .Tile_X9Y14_RAM2FAB_D2_I3(RAM2FAB_D_I[11]),
    .Tile_X9Y14_RAM2FAB_D3_I0(RAM2FAB_D_I[12]),
    .Tile_X9Y14_RAM2FAB_D3_I1(RAM2FAB_D_I[13]),
    .Tile_X9Y14_RAM2FAB_D3_I2(RAM2FAB_D_I[14]),
    .Tile_X9Y14_RAM2FAB_D3_I3(RAM2FAB_D_I[15]),
    .Tile_X9Y13_RAM2FAB_D0_I0(RAM2FAB_D_I[16]),
    .Tile_X9Y13_RAM2FAB_D0_I1(RAM2FAB_D_I[17]),
    .Tile_X9Y13_RAM2FAB_D0_I2(RAM2FAB_D_I[18]),
    .Tile_X9Y13_RAM2FAB_D0_I3(RAM2FAB_D_I[19]),
    .Tile_X9Y13_RAM2FAB_D1_I0(RAM2FAB_D_I[20]),
    .Tile_X9Y13_RAM2FAB_D1_I1(RAM2FAB_D_I[21]),
    .Tile_X9Y13_RAM2FAB_D1_I2(RAM2FAB_D_I[22]),
    .Tile_X9Y13_RAM2FAB_D1_I3(RAM2FAB_D_I[23]),
    .Tile_X9Y13_RAM2FAB_D2_I0(RAM2FAB_D_I[24]),
    .Tile_X9Y13_RAM2FAB_D2_I1(RAM2FAB_D_I[25]),
    .Tile_X9Y13_RAM2FAB_D2_I2(RAM2FAB_D_I[26]),
    .Tile_X9Y13_RAM2FAB_D2_I3(RAM2FAB_D_I[27]),
    .Tile_X9Y13_RAM2FAB_D3_I0(RAM2FAB_D_I[28]),
    .Tile_X9Y13_RAM2FAB_D3_I1(RAM2FAB_D_I[29]),
    .Tile_X9Y13_RAM2FAB_D3_I2(RAM2FAB_D_I[30]),
    .Tile_X9Y13_RAM2FAB_D3_I3(RAM2FAB_D_I[31]),
    .Tile_X9Y12_RAM2FAB_D0_I0(RAM2FAB_D_I[32]),
    .Tile_X9Y12_RAM2FAB_D0_I1(RAM2FAB_D_I[33]),
    .Tile_X9Y12_RAM2FAB_D0_I2(RAM2FAB_D_I[34]),
    .Tile_X9Y12_RAM2FAB_D0_I3(RAM2FAB_D_I[35]),
    .Tile_X9Y12_RAM2FAB_D1_I0(RAM2FAB_D_I[36]),
    .Tile_X9Y12_RAM2FAB_D1_I1(RAM2FAB_D_I[37]),
    .Tile_X9Y12_RAM2FAB_D1_I2(RAM2FAB_D_I[38]),
    .Tile_X9Y12_RAM2FAB_D1_I3(RAM2FAB_D_I[39]),
    .Tile_X9Y12_RAM2FAB_D2_I0(RAM2FAB_D_I[40]),
    .Tile_X9Y12_RAM2FAB_D2_I1(RAM2FAB_D_I[41]),
    .Tile_X9Y12_RAM2FAB_D2_I2(RAM2FAB_D_I[42]),
    .Tile_X9Y12_RAM2FAB_D2_I3(RAM2FAB_D_I[43]),
    .Tile_X9Y12_RAM2FAB_D3_I0(RAM2FAB_D_I[44]),
    .Tile_X9Y12_RAM2FAB_D3_I1(RAM2FAB_D_I[45]),
    .Tile_X9Y12_RAM2FAB_D3_I2(RAM2FAB_D_I[46]),
    .Tile_X9Y12_RAM2FAB_D3_I3(RAM2FAB_D_I[47]),
    .Tile_X9Y11_RAM2FAB_D0_I0(RAM2FAB_D_I[48]),
    .Tile_X9Y11_RAM2FAB_D0_I1(RAM2FAB_D_I[49]),
    .Tile_X9Y11_RAM2FAB_D0_I2(RAM2FAB_D_I[50]),
    .Tile_X9Y11_RAM2FAB_D0_I3(RAM2FAB_D_I[51]),
    .Tile_X9Y11_RAM2FAB_D1_I0(RAM2FAB_D_I[52]),
    .Tile_X9Y11_RAM2FAB_D1_I1(RAM2FAB_D_I[53]),
    .Tile_X9Y11_RAM2FAB_D1_I2(RAM2FAB_D_I[54]),
    .Tile_X9Y11_RAM2FAB_D1_I3(RAM2FAB_D_I[55]),
    .Tile_X9Y11_RAM2FAB_D2_I0(RAM2FAB_D_I[56]),
    .Tile_X9Y11_RAM2FAB_D2_I1(RAM2FAB_D_I[57]),
    .Tile_X9Y11_RAM2FAB_D2_I2(RAM2FAB_D_I[58]),
    .Tile_X9Y11_RAM2FAB_D2_I3(RAM2FAB_D_I[59]),
    .Tile_X9Y11_RAM2FAB_D3_I0(RAM2FAB_D_I[60]),
    .Tile_X9Y11_RAM2FAB_D3_I1(RAM2FAB_D_I[61]),
    .Tile_X9Y11_RAM2FAB_D3_I2(RAM2FAB_D_I[62]),
    .Tile_X9Y11_RAM2FAB_D3_I3(RAM2FAB_D_I[63]),
    .Tile_X9Y10_RAM2FAB_D0_I0(RAM2FAB_D_I[64]),
    .Tile_X9Y10_RAM2FAB_D0_I1(RAM2FAB_D_I[65]),
    .Tile_X9Y10_RAM2FAB_D0_I2(RAM2FAB_D_I[66]),
    .Tile_X9Y10_RAM2FAB_D0_I3(RAM2FAB_D_I[67]),
    .Tile_X9Y10_RAM2FAB_D1_I0(RAM2FAB_D_I[68]),
    .Tile_X9Y10_RAM2FAB_D1_I1(RAM2FAB_D_I[69]),
    .Tile_X9Y10_RAM2FAB_D1_I2(RAM2FAB_D_I[70]),
    .Tile_X9Y10_RAM2FAB_D1_I3(RAM2FAB_D_I[71]),
    .Tile_X9Y10_RAM2FAB_D2_I0(RAM2FAB_D_I[72]),
    .Tile_X9Y10_RAM2FAB_D2_I1(RAM2FAB_D_I[73]),
    .Tile_X9Y10_RAM2FAB_D2_I2(RAM2FAB_D_I[74]),
    .Tile_X9Y10_RAM2FAB_D2_I3(RAM2FAB_D_I[75]),
    .Tile_X9Y10_RAM2FAB_D3_I0(RAM2FAB_D_I[76]),
    .Tile_X9Y10_RAM2FAB_D3_I1(RAM2FAB_D_I[77]),
    .Tile_X9Y10_RAM2FAB_D3_I2(RAM2FAB_D_I[78]),
    .Tile_X9Y10_RAM2FAB_D3_I3(RAM2FAB_D_I[79]),
    .Tile_X9Y9_RAM2FAB_D0_I0(RAM2FAB_D_I[80]),
    .Tile_X9Y9_RAM2FAB_D0_I1(RAM2FAB_D_I[81]),
    .Tile_X9Y9_RAM2FAB_D0_I2(RAM2FAB_D_I[82]),
    .Tile_X9Y9_RAM2FAB_D0_I3(RAM2FAB_D_I[83]),
    .Tile_X9Y9_RAM2FAB_D1_I0(RAM2FAB_D_I[84]),
    .Tile_X9Y9_RAM2FAB_D1_I1(RAM2FAB_D_I[85]),
    .Tile_X9Y9_RAM2FAB_D1_I2(RAM2FAB_D_I[86]),
    .Tile_X9Y9_RAM2FAB_D1_I3(RAM2FAB_D_I[87]),
    .Tile_X9Y9_RAM2FAB_D2_I0(RAM2FAB_D_I[88]),
    .Tile_X9Y9_RAM2FAB_D2_I1(RAM2FAB_D_I[89]),
    .Tile_X9Y9_RAM2FAB_D2_I2(RAM2FAB_D_I[90]),
    .Tile_X9Y9_RAM2FAB_D2_I3(RAM2FAB_D_I[91]),
    .Tile_X9Y9_RAM2FAB_D3_I0(RAM2FAB_D_I[92]),
    .Tile_X9Y9_RAM2FAB_D3_I1(RAM2FAB_D_I[93]),
    .Tile_X9Y9_RAM2FAB_D3_I2(RAM2FAB_D_I[94]),
    .Tile_X9Y9_RAM2FAB_D3_I3(RAM2FAB_D_I[95]),
    .Tile_X9Y8_RAM2FAB_D0_I0(RAM2FAB_D_I[96]),
    .Tile_X9Y8_RAM2FAB_D0_I1(RAM2FAB_D_I[97]),
    .Tile_X9Y8_RAM2FAB_D0_I2(RAM2FAB_D_I[98]),
    .Tile_X9Y8_RAM2FAB_D0_I3(RAM2FAB_D_I[99]),
    .Tile_X9Y8_RAM2FAB_D1_I0(RAM2FAB_D_I[100]),
    .Tile_X9Y8_RAM2FAB_D1_I1(RAM2FAB_D_I[101]),
    .Tile_X9Y8_RAM2FAB_D1_I2(RAM2FAB_D_I[102]),
    .Tile_X9Y8_RAM2FAB_D1_I3(RAM2FAB_D_I[103]),
    .Tile_X9Y8_RAM2FAB_D2_I0(RAM2FAB_D_I[104]),
    .Tile_X9Y8_RAM2FAB_D2_I1(RAM2FAB_D_I[105]),
    .Tile_X9Y8_RAM2FAB_D2_I2(RAM2FAB_D_I[106]),
    .Tile_X9Y8_RAM2FAB_D2_I3(RAM2FAB_D_I[107]),
    .Tile_X9Y8_RAM2FAB_D3_I0(RAM2FAB_D_I[108]),
    .Tile_X9Y8_RAM2FAB_D3_I1(RAM2FAB_D_I[109]),
    .Tile_X9Y8_RAM2FAB_D3_I2(RAM2FAB_D_I[110]),
    .Tile_X9Y8_RAM2FAB_D3_I3(RAM2FAB_D_I[111]),
    .Tile_X9Y7_RAM2FAB_D0_I0(RAM2FAB_D_I[112]),
    .Tile_X9Y7_RAM2FAB_D0_I1(RAM2FAB_D_I[113]),
    .Tile_X9Y7_RAM2FAB_D0_I2(RAM2FAB_D_I[114]),
    .Tile_X9Y7_RAM2FAB_D0_I3(RAM2FAB_D_I[115]),
    .Tile_X9Y7_RAM2FAB_D1_I0(RAM2FAB_D_I[116]),
    .Tile_X9Y7_RAM2FAB_D1_I1(RAM2FAB_D_I[117]),
    .Tile_X9Y7_RAM2FAB_D1_I2(RAM2FAB_D_I[118]),
    .Tile_X9Y7_RAM2FAB_D1_I3(RAM2FAB_D_I[119]),
    .Tile_X9Y7_RAM2FAB_D2_I0(RAM2FAB_D_I[120]),
    .Tile_X9Y7_RAM2FAB_D2_I1(RAM2FAB_D_I[121]),
    .Tile_X9Y7_RAM2FAB_D2_I2(RAM2FAB_D_I[122]),
    .Tile_X9Y7_RAM2FAB_D2_I3(RAM2FAB_D_I[123]),
    .Tile_X9Y7_RAM2FAB_D3_I0(RAM2FAB_D_I[124]),
    .Tile_X9Y7_RAM2FAB_D3_I1(RAM2FAB_D_I[125]),
    .Tile_X9Y7_RAM2FAB_D3_I2(RAM2FAB_D_I[126]),
    .Tile_X9Y7_RAM2FAB_D3_I3(RAM2FAB_D_I[127]),
    .Tile_X9Y6_RAM2FAB_D0_I0(RAM2FAB_D_I[128]),
    .Tile_X9Y6_RAM2FAB_D0_I1(RAM2FAB_D_I[129]),
    .Tile_X9Y6_RAM2FAB_D0_I2(RAM2FAB_D_I[130]),
    .Tile_X9Y6_RAM2FAB_D0_I3(RAM2FAB_D_I[131]),
    .Tile_X9Y6_RAM2FAB_D1_I0(RAM2FAB_D_I[132]),
    .Tile_X9Y6_RAM2FAB_D1_I1(RAM2FAB_D_I[133]),
    .Tile_X9Y6_RAM2FAB_D1_I2(RAM2FAB_D_I[134]),
    .Tile_X9Y6_RAM2FAB_D1_I3(RAM2FAB_D_I[135]),
    .Tile_X9Y6_RAM2FAB_D2_I0(RAM2FAB_D_I[136]),
    .Tile_X9Y6_RAM2FAB_D2_I1(RAM2FAB_D_I[137]),
    .Tile_X9Y6_RAM2FAB_D2_I2(RAM2FAB_D_I[138]),
    .Tile_X9Y6_RAM2FAB_D2_I3(RAM2FAB_D_I[139]),
    .Tile_X9Y6_RAM2FAB_D3_I0(RAM2FAB_D_I[140]),
    .Tile_X9Y6_RAM2FAB_D3_I1(RAM2FAB_D_I[141]),
    .Tile_X9Y6_RAM2FAB_D3_I2(RAM2FAB_D_I[142]),
    .Tile_X9Y6_RAM2FAB_D3_I3(RAM2FAB_D_I[143]),
    .Tile_X9Y5_RAM2FAB_D0_I0(RAM2FAB_D_I[144]),
    .Tile_X9Y5_RAM2FAB_D0_I1(RAM2FAB_D_I[145]),
    .Tile_X9Y5_RAM2FAB_D0_I2(RAM2FAB_D_I[146]),
    .Tile_X9Y5_RAM2FAB_D0_I3(RAM2FAB_D_I[147]),
    .Tile_X9Y5_RAM2FAB_D1_I0(RAM2FAB_D_I[148]),
    .Tile_X9Y5_RAM2FAB_D1_I1(RAM2FAB_D_I[149]),
    .Tile_X9Y5_RAM2FAB_D1_I2(RAM2FAB_D_I[150]),
    .Tile_X9Y5_RAM2FAB_D1_I3(RAM2FAB_D_I[151]),
    .Tile_X9Y5_RAM2FAB_D2_I0(RAM2FAB_D_I[152]),
    .Tile_X9Y5_RAM2FAB_D2_I1(RAM2FAB_D_I[153]),
    .Tile_X9Y5_RAM2FAB_D2_I2(RAM2FAB_D_I[154]),
    .Tile_X9Y5_RAM2FAB_D2_I3(RAM2FAB_D_I[155]),
    .Tile_X9Y5_RAM2FAB_D3_I0(RAM2FAB_D_I[156]),
    .Tile_X9Y5_RAM2FAB_D3_I1(RAM2FAB_D_I[157]),
    .Tile_X9Y5_RAM2FAB_D3_I2(RAM2FAB_D_I[158]),
    .Tile_X9Y5_RAM2FAB_D3_I3(RAM2FAB_D_I[159]),
    .Tile_X9Y4_RAM2FAB_D0_I0(RAM2FAB_D_I[160]),
    .Tile_X9Y4_RAM2FAB_D0_I1(RAM2FAB_D_I[161]),
    .Tile_X9Y4_RAM2FAB_D0_I2(RAM2FAB_D_I[162]),
    .Tile_X9Y4_RAM2FAB_D0_I3(RAM2FAB_D_I[163]),
    .Tile_X9Y4_RAM2FAB_D1_I0(RAM2FAB_D_I[164]),
    .Tile_X9Y4_RAM2FAB_D1_I1(RAM2FAB_D_I[165]),
    .Tile_X9Y4_RAM2FAB_D1_I2(RAM2FAB_D_I[166]),
    .Tile_X9Y4_RAM2FAB_D1_I3(RAM2FAB_D_I[167]),
    .Tile_X9Y4_RAM2FAB_D2_I0(RAM2FAB_D_I[168]),
    .Tile_X9Y4_RAM2FAB_D2_I1(RAM2FAB_D_I[169]),
    .Tile_X9Y4_RAM2FAB_D2_I2(RAM2FAB_D_I[170]),
    .Tile_X9Y4_RAM2FAB_D2_I3(RAM2FAB_D_I[171]),
    .Tile_X9Y4_RAM2FAB_D3_I0(RAM2FAB_D_I[172]),
    .Tile_X9Y4_RAM2FAB_D3_I1(RAM2FAB_D_I[173]),
    .Tile_X9Y4_RAM2FAB_D3_I2(RAM2FAB_D_I[174]),
    .Tile_X9Y4_RAM2FAB_D3_I3(RAM2FAB_D_I[175]),
    .Tile_X9Y3_RAM2FAB_D0_I0(RAM2FAB_D_I[176]),
    .Tile_X9Y3_RAM2FAB_D0_I1(RAM2FAB_D_I[177]),
    .Tile_X9Y3_RAM2FAB_D0_I2(RAM2FAB_D_I[178]),
    .Tile_X9Y3_RAM2FAB_D0_I3(RAM2FAB_D_I[179]),
    .Tile_X9Y3_RAM2FAB_D1_I0(RAM2FAB_D_I[180]),
    .Tile_X9Y3_RAM2FAB_D1_I1(RAM2FAB_D_I[181]),
    .Tile_X9Y3_RAM2FAB_D1_I2(RAM2FAB_D_I[182]),
    .Tile_X9Y3_RAM2FAB_D1_I3(RAM2FAB_D_I[183]),
    .Tile_X9Y3_RAM2FAB_D2_I0(RAM2FAB_D_I[184]),
    .Tile_X9Y3_RAM2FAB_D2_I1(RAM2FAB_D_I[185]),
    .Tile_X9Y3_RAM2FAB_D2_I2(RAM2FAB_D_I[186]),
    .Tile_X9Y3_RAM2FAB_D2_I3(RAM2FAB_D_I[187]),
    .Tile_X9Y3_RAM2FAB_D3_I0(RAM2FAB_D_I[188]),
    .Tile_X9Y3_RAM2FAB_D3_I1(RAM2FAB_D_I[189]),
    .Tile_X9Y3_RAM2FAB_D3_I2(RAM2FAB_D_I[190]),
    .Tile_X9Y3_RAM2FAB_D3_I3(RAM2FAB_D_I[191]),
    .Tile_X9Y2_RAM2FAB_D0_I0(RAM2FAB_D_I[192]),
    .Tile_X9Y2_RAM2FAB_D0_I1(RAM2FAB_D_I[193]),
    .Tile_X9Y2_RAM2FAB_D0_I2(RAM2FAB_D_I[194]),
    .Tile_X9Y2_RAM2FAB_D0_I3(RAM2FAB_D_I[195]),
    .Tile_X9Y2_RAM2FAB_D1_I0(RAM2FAB_D_I[196]),
    .Tile_X9Y2_RAM2FAB_D1_I1(RAM2FAB_D_I[197]),
    .Tile_X9Y2_RAM2FAB_D1_I2(RAM2FAB_D_I[198]),
    .Tile_X9Y2_RAM2FAB_D1_I3(RAM2FAB_D_I[199]),
    .Tile_X9Y2_RAM2FAB_D2_I0(RAM2FAB_D_I[200]),
    .Tile_X9Y2_RAM2FAB_D2_I1(RAM2FAB_D_I[201]),
    .Tile_X9Y2_RAM2FAB_D2_I2(RAM2FAB_D_I[202]),
    .Tile_X9Y2_RAM2FAB_D2_I3(RAM2FAB_D_I[203]),
    .Tile_X9Y2_RAM2FAB_D3_I0(RAM2FAB_D_I[204]),
    .Tile_X9Y2_RAM2FAB_D3_I1(RAM2FAB_D_I[205]),
    .Tile_X9Y2_RAM2FAB_D3_I2(RAM2FAB_D_I[206]),
    .Tile_X9Y2_RAM2FAB_D3_I3(RAM2FAB_D_I[207]),
    .Tile_X9Y1_RAM2FAB_D0_I0(RAM2FAB_D_I[208]),
    .Tile_X9Y1_RAM2FAB_D0_I1(RAM2FAB_D_I[209]),
    .Tile_X9Y1_RAM2FAB_D0_I2(RAM2FAB_D_I[210]),
    .Tile_X9Y1_RAM2FAB_D0_I3(RAM2FAB_D_I[211]),
    .Tile_X9Y1_RAM2FAB_D1_I0(RAM2FAB_D_I[212]),
    .Tile_X9Y1_RAM2FAB_D1_I1(RAM2FAB_D_I[213]),
    .Tile_X9Y1_RAM2FAB_D1_I2(RAM2FAB_D_I[214]),
    .Tile_X9Y1_RAM2FAB_D1_I3(RAM2FAB_D_I[215]),
    .Tile_X9Y1_RAM2FAB_D2_I0(RAM2FAB_D_I[216]),
    .Tile_X9Y1_RAM2FAB_D2_I1(RAM2FAB_D_I[217]),
    .Tile_X9Y1_RAM2FAB_D2_I2(RAM2FAB_D_I[218]),
    .Tile_X9Y1_RAM2FAB_D2_I3(RAM2FAB_D_I[219]),
    .Tile_X9Y1_RAM2FAB_D3_I0(RAM2FAB_D_I[220]),
    .Tile_X9Y1_RAM2FAB_D3_I1(RAM2FAB_D_I[221]),
    .Tile_X9Y1_RAM2FAB_D3_I2(RAM2FAB_D_I[222]),
    .Tile_X9Y1_RAM2FAB_D3_I3(RAM2FAB_D_I[223]),
    .Tile_X0Y14_B_T_top(T_top[0]),
    .Tile_X0Y14_A_T_top(T_top[1]),
    .Tile_X0Y13_B_T_top(T_top[2]),
    .Tile_X0Y13_A_T_top(T_top[3]),
    .Tile_X0Y12_B_T_top(T_top[4]),
    .Tile_X0Y12_A_T_top(T_top[5]),
    .Tile_X0Y11_B_T_top(T_top[6]),
    .Tile_X0Y11_A_T_top(T_top[7]),
    .Tile_X0Y10_B_T_top(T_top[8]),
    .Tile_X0Y10_A_T_top(T_top[9]),
    .Tile_X0Y9_B_T_top(T_top[10]),
    .Tile_X0Y9_A_T_top(T_top[11]),
    .Tile_X0Y8_B_T_top(T_top[12]),
    .Tile_X0Y8_A_T_top(T_top[13]),
    .Tile_X0Y7_B_T_top(T_top[14]),
    .Tile_X0Y7_A_T_top(T_top[15]),
    .Tile_X0Y6_B_T_top(T_top[16]),
    .Tile_X0Y6_A_T_top(T_top[17]),
    .Tile_X0Y5_B_T_top(T_top[18]),
    .Tile_X0Y5_A_T_top(T_top[19]),
    .Tile_X0Y4_B_T_top(T_top[20]),
    .Tile_X0Y4_A_T_top(T_top[21]),
    .Tile_X0Y3_B_T_top(T_top[22]),
    .Tile_X0Y3_A_T_top(T_top[23]),
    .Tile_X0Y2_B_T_top(T_top[24]),
    .Tile_X0Y2_A_T_top(T_top[25]),
    .Tile_X0Y1_B_T_top(T_top[26]),
    .Tile_X0Y1_A_T_top(T_top[27]),
    .UserCLK(CLK),
    .FrameData(FrameData),
    .FrameStrobe(FrameSelect)
);


BlockRAM_1KB Inst_BlockRAM_0 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[7:0]),
    .rd_data(RAM2FAB_D_I[31:0]),
    .wr_addr(FAB2RAM_A_O[15:8]),
    .wr_data(FAB2RAM_D_O[31:0]),
    .C0(FAB2RAM_C_O[0]),
    .C1(FAB2RAM_C_O[1]),
    .C2(FAB2RAM_C_O[2]),
    .C3(FAB2RAM_C_O[3]),
    .C4(FAB2RAM_C_O[4]),
    .C5(FAB2RAM_C_O[5])
);

BlockRAM_1KB Inst_BlockRAM_1 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[23:16]),
    .rd_data(RAM2FAB_D_I[63:32]),
    .wr_addr(FAB2RAM_A_O[31:24]),
    .wr_data(FAB2RAM_D_O[63:32]),
    .C0(FAB2RAM_C_O[8]),
    .C1(FAB2RAM_C_O[9]),
    .C2(FAB2RAM_C_O[10]),
    .C3(FAB2RAM_C_O[11]),
    .C4(FAB2RAM_C_O[12]),
    .C5(FAB2RAM_C_O[13])
);

BlockRAM_1KB Inst_BlockRAM_2 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[39:32]),
    .rd_data(RAM2FAB_D_I[95:64]),
    .wr_addr(FAB2RAM_A_O[47:40]),
    .wr_data(FAB2RAM_D_O[95:64]),
    .C0(FAB2RAM_C_O[16]),
    .C1(FAB2RAM_C_O[17]),
    .C2(FAB2RAM_C_O[18]),
    .C3(FAB2RAM_C_O[19]),
    .C4(FAB2RAM_C_O[20]),
    .C5(FAB2RAM_C_O[21])
);

BlockRAM_1KB Inst_BlockRAM_3 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[55:48]),
    .rd_data(RAM2FAB_D_I[127:96]),
    .wr_addr(FAB2RAM_A_O[63:56]),
    .wr_data(FAB2RAM_D_O[127:96]),
    .C0(FAB2RAM_C_O[24]),
    .C1(FAB2RAM_C_O[25]),
    .C2(FAB2RAM_C_O[26]),
    .C3(FAB2RAM_C_O[27]),
    .C4(FAB2RAM_C_O[28]),
    .C5(FAB2RAM_C_O[29])
);

BlockRAM_1KB Inst_BlockRAM_4 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[71:64]),
    .rd_data(RAM2FAB_D_I[159:128]),
    .wr_addr(FAB2RAM_A_O[79:72]),
    .wr_data(FAB2RAM_D_O[159:128]),
    .C0(FAB2RAM_C_O[32]),
    .C1(FAB2RAM_C_O[33]),
    .C2(FAB2RAM_C_O[34]),
    .C3(FAB2RAM_C_O[35]),
    .C4(FAB2RAM_C_O[36]),
    .C5(FAB2RAM_C_O[37])
);

BlockRAM_1KB Inst_BlockRAM_5 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[87:80]),
    .rd_data(RAM2FAB_D_I[191:160]),
    .wr_addr(FAB2RAM_A_O[95:88]),
    .wr_data(FAB2RAM_D_O[191:160]),
    .C0(FAB2RAM_C_O[40]),
    .C1(FAB2RAM_C_O[41]),
    .C2(FAB2RAM_C_O[42]),
    .C3(FAB2RAM_C_O[43]),
    .C4(FAB2RAM_C_O[44]),
    .C5(FAB2RAM_C_O[45])
);

BlockRAM_1KB Inst_BlockRAM_6 (
    .clk(CLK),
    .rd_addr(FAB2RAM_A_O[103:96]),
    .rd_data(RAM2FAB_D_I[223:192]),
    .wr_addr(FAB2RAM_A_O[111:104]),
    .wr_data(FAB2RAM_D_O[223:192]),
    .C0(FAB2RAM_C_O[48]),
    .C1(FAB2RAM_C_O[49]),
    .C2(FAB2RAM_C_O[50]),
    .C3(FAB2RAM_C_O[51]),
    .C4(FAB2RAM_C_O[52]),
    .C5(FAB2RAM_C_O[53])
);

assign FrameData = {32'h12345678,FrameRegister,32'h12345678};
endmodule