module S_IO_switch_matrix #(
    parameter NoConfigBits = 0
)(

);

localparam reg GND0 = 0;
localparam reg GND = 0;
localparam reg VCC0 = 1;
localparam reg VCC = 1;
localparam reg VDD0 = 1;
localparam reg VDD = 1;

endmodule
