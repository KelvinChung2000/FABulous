(* blackbox *)
module reg_unit #(
)
(
    input en,
    input [31:0] reg_in,
    input rst,
    output [31:0] reg_out,
    input clk
);

endmodule
