module accumulate #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] i3_add;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i4_data_size1;
wire[WIDTH-1:0] i4_mul1;
wire[WIDTH-1:0] i4_add1;
wire[WIDTH-1:0] i5_load;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i6_add;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i7_data_size1;
wire[WIDTH-1:0] i7_mul1;
wire[WIDTH-1:0] i7_add1;
wire[WIDTH-1:0] i8_load;
wire[WIDTH-1:0] i9_add;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i10_data_size1;
wire[WIDTH-1:0] i10_mul1;
wire[WIDTH-1:0] i10_add1;
wire[WIDTH-1:0] i11_load;
wire[WIDTH-1:0] i12_mul;
wire[WIDTH-1:0] i14_add;
wire[WIDTH-1:0] input0;
wire i15_icmp;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] i3_add_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i4_data_size1_alu;
wire[WIDTH-1:0] i4_mul1_alu;
wire[WIDTH-1:0] i4_add1_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i6_add_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i7_data_size1_alu;
wire[WIDTH-1:0] i7_mul1_alu;
wire[WIDTH-1:0] i7_add1_alu;
wire[WIDTH-1:0] i9_add_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i10_data_size1_alu;
wire[WIDTH-1:0] i10_mul1_alu;
wire[WIDTH-1:0] i10_add1_alu;
wire[WIDTH-1:0] i12_mul_alu;
wire[WIDTH-1:0] i14_add_alu;
wire[WIDTH-1:0] i14_output_alu;
wire[WIDTH-1:0] i13_store;
wire[WIDTH-1:0] i16_br;
wire[WIDTH-1:0] i14_output;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(1)) inst_const0(.const_out(const0));
ALU #(.ALU_func(add_op)) inst_i3_add(.data_in1(const0), .data_in2(i3_add), .data_in3(), .data_out(i3_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add_reg(.reg_in(i3_add_alu), .reg_out(i3_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2560)) inst_const2(.const_out(const2));
const_unit #(.ConfigBits(4)) inst_i4_data_size1(.const_out(i4_data_size1));
ALU #(.ALU_func(mul_op)) inst_i4_mul1(.data_in1(i3_add), .data_in2(i4_data_size1), .data_in3(), .data_out(i4_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_mul1_reg(.reg_in(i4_mul1_alu), .reg_out(i4_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i4_add1(.data_in1(const2), .data_in2(i4_mul1), .data_in3(), .data_out(i4_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_add1_reg(.reg_in(i4_add1_alu), .reg_out(i4_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i5_load(.addr0(i4_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i5_load));
const_unit #(.ConfigBits(0)) inst_const3(.const_out(const3));
ALU #(.ALU_func(add_op)) inst_i6_add(.data_in1(const3), .data_in2(i3_add), .data_in3(), .data_out(i6_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add_reg(.reg_in(i6_add_alu), .reg_out(i6_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2816)) inst_const4(.const_out(const4));
const_unit #(.ConfigBits(4)) inst_i7_data_size1(.const_out(i7_data_size1));
ALU #(.ALU_func(mul_op)) inst_i7_mul1(.data_in1(i6_add), .data_in2(i7_data_size1), .data_in3(), .data_out(i7_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_mul1_reg(.reg_in(i7_mul1_alu), .reg_out(i7_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i7_add1(.data_in1(const4), .data_in2(i7_mul1), .data_in3(), .data_out(i7_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i7_add1_reg(.reg_in(i7_add1_alu), .reg_out(i7_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i8_load(.addr0(i7_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i8_load));
ALU #(.ALU_func(add_op)) inst_i9_add(.data_in1(i5_load), .data_in2(i8_load), .data_in3(), .data_out(i9_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add_reg(.reg_in(i9_add_alu), .reg_out(i9_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(3072)) inst_const5(.const_out(const5));
const_unit #(.ConfigBits(4)) inst_i10_data_size1(.const_out(i10_data_size1));
ALU #(.ALU_func(mul_op)) inst_i10_mul1(.data_in1(i10_data_size1), .data_in2(i3_add), .data_in3(), .data_out(i10_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_mul1_reg(.reg_in(i10_mul1_alu), .reg_out(i10_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i10_add1(.data_in1(const5), .data_in2(i10_mul1), .data_in3(), .data_out(i10_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_add1_reg(.reg_in(i10_add1_alu), .reg_out(i10_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i11_load(.addr0(i10_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i11_load));
ALU #(.ALU_func(mul_op)) inst_i12_mul(.data_in1(i9_add), .data_in2(i11_load), .data_in3(), .data_out(i12_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_mul_reg(.reg_in(i12_mul_alu), .reg_out(i12_mul), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i13_store(.addr0(i10_add1), .reset(global_rst), .write_data(i12_mul), .write_en(), .read_data(i13_store));
ALU #(.ALU_func(add_op)) inst_i14_add(.data_in1(i12_mul), .data_in2(i14_add), .data_in3(), .data_out(i14_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_add_reg(.reg_in(i14_add_alu), .reg_out(i14_add), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i15_icmp(.A(i3_add), .B(input0), .Y(i15_icmp));
(* keep *) IO_WIDTH_1 inst_i16_br(.from_fabric(i15_icmp), .in(), .to_fabric(), .out());
(* keep *) IO inst_i14_output(.from_fabric(i14_add), .in(), .to_fabric(), .out());

endmodule
