module conv3 #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const1;
wire[WIDTH-1:0] i2_data_size1;
wire[WIDTH-1:0] i2_mul1;
wire[WIDTH-1:0] i2_add1;
wire[WIDTH-1:0] i3_load;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i4_mul;
wire[WIDTH-1:0] i5_add;
wire[WIDTH-1:0] i6_data_size1;
wire[WIDTH-1:0] i6_mul1;
wire[WIDTH-1:0] i6_add1;
wire[WIDTH-1:0] i7_load;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i8_mul;
wire[WIDTH-1:0] i9_add;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i10_add;
wire[WIDTH-1:0] i11_data_size1;
wire[WIDTH-1:0] i11_mul1;
wire[WIDTH-1:0] i11_add1;
wire[WIDTH-1:0] i12_load;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i13_mul;
wire[WIDTH-1:0] i14_add;
wire[WIDTH-1:0] const6;
wire[WIDTH-1:0] i15_data_size1;
wire[WIDTH-1:0] i15_mul1;
wire[WIDTH-1:0] i15_add1;
wire[WIDTH-1:0] input0;
wire i17_icmp;
wire[WIDTH-1:0] const1_dup_1;
wire[WIDTH-1:0] const1_dup_2;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const1_alu;
wire[WIDTH-1:0] i2_data_size1_alu;
wire[WIDTH-1:0] i2_mul1_alu;
wire[WIDTH-1:0] i2_add1_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i4_mul_alu;
wire[WIDTH-1:0] i5_add_alu;
wire[WIDTH-1:0] i6_data_size1_alu;
wire[WIDTH-1:0] i6_mul1_alu;
wire[WIDTH-1:0] i6_add1_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i8_mul_alu;
wire[WIDTH-1:0] i9_add_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i10_add_alu;
wire[WIDTH-1:0] i11_data_size1_alu;
wire[WIDTH-1:0] i11_mul1_alu;
wire[WIDTH-1:0] i11_add1_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i13_mul_alu;
wire[WIDTH-1:0] i14_add_alu;
wire[WIDTH-1:0] const6_alu;
wire[WIDTH-1:0] i15_data_size1_alu;
wire[WIDTH-1:0] i15_mul1_alu;
wire[WIDTH-1:0] i15_add1_alu;
wire[WIDTH-1:0] const1_dup_1_alu;
wire[WIDTH-1:0] const1_dup_2_alu;
wire[WIDTH-1:0] i16_store;
wire[WIDTH-1:0] i18_br;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(1)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const1(.const_out(const1));
const_unit #(.ConfigBits(4)) inst_i2_data_size1(.const_out(i2_data_size1));
ALU #(.ALU_func(mul_op)) inst_i2_mul1(.data_in1(i2_data_size1), .data_in2(i5_add), .data_in3(), .data_out(i2_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i2_mul1_reg(.reg_in(i2_mul1_alu), .reg_out(i2_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i2_add1(.data_in1(const1), .data_in2(i2_mul1), .data_in3(), .data_out(i2_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i2_add1_reg(.reg_in(i2_add1_alu), .reg_out(i2_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i3_load(.addr0(i2_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i3_load));
const_unit #(.ConfigBits(10)) inst_const2(.const_out(const2));
ALU #(.ALU_func(mul_op)) inst_i4_mul(.data_in1(i3_load), .data_in2(const2), .data_in3(), .data_out(i4_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_mul_reg(.reg_in(i4_mul_alu), .reg_out(i4_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i5_add(.data_in1(const0), .data_in2(i5_add), .data_in3(), .data_out(i5_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_add_reg(.reg_in(i5_add_alu), .reg_out(i5_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i6_data_size1(.const_out(i6_data_size1));
ALU #(.ALU_func(mul_op)) inst_i6_mul1(.data_in1(i5_add), .data_in2(i6_data_size1), .data_in3(), .data_out(i6_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_mul1_reg(.reg_in(i6_mul1_alu), .reg_out(i6_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i6_add1(.data_in1(i6_mul1), .data_in2(const1_dup_1), .data_in3(), .data_out(i6_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add1_reg(.reg_in(i6_add1_alu), .reg_out(i6_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i7_load(.addr0(i6_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i7_load));
const_unit #(.ConfigBits(20)) inst_const3(.const_out(const3));
ALU #(.ALU_func(mul_op)) inst_i8_mul(.data_in1(i7_load), .data_in2(const3), .data_in3(), .data_out(i8_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_mul_reg(.reg_in(i8_mul_alu), .reg_out(i8_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i9_add(.data_in1(i4_mul), .data_in2(i8_mul), .data_in3(), .data_out(i9_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add_reg(.reg_in(i9_add_alu), .reg_out(i9_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2)) inst_const4(.const_out(const4));
ALU #(.ALU_func(add_op)) inst_i10_add(.data_in1(const4), .data_in2(i5_add), .data_in3(), .data_out(i10_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_add_reg(.reg_in(i10_add_alu), .reg_out(i10_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i11_data_size1(.const_out(i11_data_size1));
ALU #(.ALU_func(mul_op)) inst_i11_mul1(.data_in1(i10_add), .data_in2(i11_data_size1), .data_in3(), .data_out(i11_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_mul1_reg(.reg_in(i11_mul1_alu), .reg_out(i11_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i11_add1(.data_in1(i11_mul1), .data_in2(const1_dup_2), .data_in3(), .data_out(i11_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_add1_reg(.reg_in(i11_add1_alu), .reg_out(i11_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i12_load(.addr0(i11_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i12_load));
const_unit #(.ConfigBits(3)) inst_const5(.const_out(const5));
ALU #(.ALU_func(mul_op)) inst_i13_mul(.data_in1(i12_load), .data_in2(const5), .data_in3(), .data_out(i13_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i13_mul_reg(.reg_in(i13_mul_alu), .reg_out(i13_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i14_add(.data_in1(i9_add), .data_in2(i13_mul), .data_in3(), .data_out(i14_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_add_reg(.reg_in(i14_add_alu), .reg_out(i14_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2816)) inst_const6(.const_out(const6));
const_unit #(.ConfigBits(4)) inst_i15_data_size1(.const_out(i15_data_size1));
ALU #(.ALU_func(mul_op)) inst_i15_mul1(.data_in1(i15_data_size1), .data_in2(i5_add), .data_in3(), .data_out(i15_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_mul1_reg(.reg_in(i15_mul1_alu), .reg_out(i15_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i15_add1(.data_in1(const6), .data_in2(i15_mul1), .data_in3(), .data_out(i15_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_add1_reg(.reg_in(i15_add1_alu), .reg_out(i15_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i16_store(.addr0(i14_add), .reset(global_rst), .write_data(i15_add1), .write_en(), .read_data(i16_store));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i17_icmp(.A(i5_add), .B(input0), .Y(i17_icmp));
(* keep *) IO_WIDTH_1 inst_i18_br(.from_fabric(i17_icmp), .in(), .to_fabric(), .out());
const_unit #(.ConfigBits(2560)) inst_const1_dup_1(.const_out(const1_dup_1));
const_unit #(.ConfigBits(2560)) inst_const1_dup_2(.const_out(const1_dup_2));

endmodule
