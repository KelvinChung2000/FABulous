(* blackbox *)
module Mem #(
    parameter config_bits = 0
)
(
    input wire[31:0] addr0,
    input wire reset,
    input wire[31:0] write_data,
    input wire write_en,
    output reg[31:0] read_data
);

endmodule


(* blackbox *)
module IO #(
)
(
    input wire[31:0] from_fabric,
    input wire[31:0] in,
    output reg[31:0] to_fabric,
    output reg[31:0] out
);

endmodule


(* blackbox *)
module IO_WIDTH_1 #(
)
(
    input wire from_fabric,
    input wire in,
    output reg to_fabric,
    output reg out
);

endmodule


(* blackbox *)
module ALU #(
    parameter ALU_func = 0
)
(
    input wire[31:0] data_in1,
    input wire[31:0] data_in2,
    input wire data_in3,
    output reg[31:0] data_out
);

endmodule


(* blackbox *)
module compare #(
    parameter conf = 0
)
(
    input wire[31:0] A,
    input wire[31:0] B,
    output reg Y
);

endmodule


(* blackbox *)
module const_unit #(
    parameter ConfigBits = 0
)
(
    output reg[31:0] const_out
);

endmodule


(* blackbox *)
module logic_op #(
    parameter conf = 0
)
(
    input wire A,
    input wire B,
    output reg Y
);

endmodule


(* blackbox *)
module reg_unit #(
    parameter tide_en = 0,
    parameter tide_rst = 0
)
(
    input wire[31:0] reg_in,
    output reg[31:0] reg_out,
    input wire en,
    input wire rst
);

endmodule


(* blackbox *)
module reg_unit_WIDTH_1 #(
    parameter tide_en = 0,
    parameter tide_rst = 0
)
(
    input wire reg_in,
    output reg reg_out,
    input wire en,
    input wire rst
);

endmodule


