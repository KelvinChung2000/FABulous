module mac2 #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i4_data_size1;
wire[WIDTH-1:0] i4_mul1;
wire[WIDTH-1:0] i4_add1;
wire[WIDTH-1:0] i5_load;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i6_data_size1;
wire[WIDTH-1:0] i6_mul1;
wire[WIDTH-1:0] i6_add1;
wire[WIDTH-1:0] i7_load;
wire[WIDTH-1:0] i8_mul;
wire[WIDTH-1:0] i9_add;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i10_add;
wire[WIDTH-1:0] i11_mul;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i12_data_size1;
wire[WIDTH-1:0] i12_mul1;
wire[WIDTH-1:0] i12_add1;
wire[WIDTH-1:0] i13_load;
wire[WIDTH-1:0] i14_mul;
wire[WIDTH-1:0] const6;
wire[WIDTH-1:0] i15_data_size1;
wire[WIDTH-1:0] i15_mul1;
wire[WIDTH-1:0] i15_add1;
wire[WIDTH-1:0] i16_load;
wire[WIDTH-1:0] i17_mul;
wire[WIDTH-1:0] i18_add;
wire[WIDTH-1:0] i19_add;
wire[WIDTH-1:0] input0;
wire i20_icmp;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i4_data_size1_alu;
wire[WIDTH-1:0] i4_mul1_alu;
wire[WIDTH-1:0] i4_add1_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i6_data_size1_alu;
wire[WIDTH-1:0] i6_mul1_alu;
wire[WIDTH-1:0] i6_add1_alu;
wire[WIDTH-1:0] i8_mul_alu;
wire[WIDTH-1:0] i9_add_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i10_add_alu;
wire[WIDTH-1:0] i11_mul_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i12_data_size1_alu;
wire[WIDTH-1:0] i12_mul1_alu;
wire[WIDTH-1:0] i12_add1_alu;
wire[WIDTH-1:0] i14_mul_alu;
wire[WIDTH-1:0] const6_alu;
wire[WIDTH-1:0] i15_data_size1_alu;
wire[WIDTH-1:0] i15_mul1_alu;
wire[WIDTH-1:0] i15_add1_alu;
wire[WIDTH-1:0] i17_mul_alu;
wire[WIDTH-1:0] i18_add_alu;
wire[WIDTH-1:0] i19_add_alu;
wire[WIDTH-1:0] i9_output_alu;
wire[WIDTH-1:0] i18_output_alu;
wire[WIDTH-1:0] i21_br;
wire[WIDTH-1:0] i9_output;
wire[WIDTH-1:0] i18_output;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(1)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const2(.const_out(const2));
const_unit #(.ConfigBits(4)) inst_i4_data_size1(.const_out(i4_data_size1));
ALU #(.ALU_func(mul_op)) inst_i4_mul1(.data_in1(i4_data_size1), .data_in2(i19_add), .data_in3(), .data_out(i4_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_mul1_reg(.reg_in(i4_mul1_alu), .reg_out(i4_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i4_add1(.data_in1(const2), .data_in2(i4_mul1), .data_in3(), .data_out(i4_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i4_add1_reg(.reg_in(i4_add1_alu), .reg_out(i4_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i5_load(.addr0(i4_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i5_load));
const_unit #(.ConfigBits(2816)) inst_const3(.const_out(const3));
const_unit #(.ConfigBits(4)) inst_i6_data_size1(.const_out(i6_data_size1));
ALU #(.ALU_func(mul_op)) inst_i6_mul1(.data_in1(i6_data_size1), .data_in2(i19_add), .data_in3(), .data_out(i6_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_mul1_reg(.reg_in(i6_mul1_alu), .reg_out(i6_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i6_add1(.data_in1(const3), .data_in2(i6_mul1), .data_in3(), .data_out(i6_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add1_reg(.reg_in(i6_add1_alu), .reg_out(i6_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i7_load(.addr0(i6_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i7_load));
ALU #(.ALU_func(mul_op)) inst_i8_mul(.data_in1(i5_load), .data_in2(i7_load), .data_in3(), .data_out(i8_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_mul_reg(.reg_in(i8_mul_alu), .reg_out(i8_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i9_add(.data_in1(i8_mul), .data_in2(i9_add), .data_in3(), .data_out(i9_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add_reg(.reg_in(i9_add_alu), .reg_out(i9_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(1)) inst_const4(.const_out(const4));
ALU #(.ALU_func(add_op)) inst_i10_add(.data_in1(i7_load), .data_in2(const4), .data_in3(), .data_out(i10_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i10_add_reg(.reg_in(i10_add_alu), .reg_out(i10_add), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i11_mul(.data_in1(i5_load), .data_in2(i10_add), .data_in3(), .data_out(i11_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_mul_reg(.reg_in(i11_mul_alu), .reg_out(i11_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(3072)) inst_const5(.const_out(const5));
const_unit #(.ConfigBits(4)) inst_i12_data_size1(.const_out(i12_data_size1));
ALU #(.ALU_func(mul_op)) inst_i12_mul1(.data_in1(i12_data_size1), .data_in2(i19_add), .data_in3(), .data_out(i12_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_mul1_reg(.reg_in(i12_mul1_alu), .reg_out(i12_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i12_add1(.data_in1(const5), .data_in2(i12_mul1), .data_in3(), .data_out(i12_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_add1_reg(.reg_in(i12_add1_alu), .reg_out(i12_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i13_load(.addr0(i12_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i13_load));
ALU #(.ALU_func(mul_op)) inst_i14_mul(.data_in1(i11_mul), .data_in2(i13_load), .data_in3(), .data_out(i14_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_mul_reg(.reg_in(i14_mul_alu), .reg_out(i14_mul), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(3328)) inst_const6(.const_out(const6));
const_unit #(.ConfigBits(4)) inst_i15_data_size1(.const_out(i15_data_size1));
ALU #(.ALU_func(mul_op)) inst_i15_mul1(.data_in1(i15_data_size1), .data_in2(i19_add), .data_in3(), .data_out(i15_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_mul1_reg(.reg_in(i15_mul1_alu), .reg_out(i15_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i15_add1(.data_in1(const6), .data_in2(i15_mul1), .data_in3(), .data_out(i15_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_add1_reg(.reg_in(i15_add1_alu), .reg_out(i15_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i16_load(.addr0(i15_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i16_load));
ALU #(.ALU_func(mul_op)) inst_i17_mul(.data_in1(i14_mul), .data_in2(i16_load), .data_in3(), .data_out(i17_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i17_mul_reg(.reg_in(i17_mul_alu), .reg_out(i17_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i18_add(.data_in1(i17_mul), .data_in2(i18_add), .data_in3(), .data_out(i18_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i18_add_reg(.reg_in(i18_add_alu), .reg_out(i18_add), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i19_add(.data_in1(const0), .data_in2(i19_add), .data_in3(), .data_out(i19_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i19_add_reg(.reg_in(i19_add_alu), .reg_out(i19_add), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i20_icmp(.A(i19_add), .B(input0), .Y(i20_icmp));
(* keep *) IO_WIDTH_1 inst_i21_br(.from_fabric(i20_icmp), .in(), .to_fabric(), .out());
(* keep *) IO inst_i9_output(.from_fabric(i9_add), .in(), .to_fabric(), .out());
(* keep *) IO inst_i18_output(.from_fabric(i18_add), .in(), .to_fabric(), .out());

endmodule
