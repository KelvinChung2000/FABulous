module hycube_wrapper #(
    parameter include_eFPGA = 1,
    parameter NumberOfCols = 6,
    parameter NumberOfRows = 6,
    parameter FrameBitsPerRow = 32,
    parameter MaxFramePerCol = 32,
    parameter FrameSelectWidth = 6,
    parameter RowSelectWidth = 3,
    parameter desync_flag = 20
)(

);


endmodule
