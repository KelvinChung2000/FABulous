module mults2 #(parameter WIDTH=32);

localparam add_op = 0;
localparam const_op = 1;
localparam icmp_op = 2;
localparam io_width_1_op = 3;
localparam mul_op = 4;

wire global_en;
wire global_rst;

wire[WIDTH-1:0] const0;
wire[WIDTH-1:0] const2;
wire[WIDTH-1:0] i3_data_size1;
wire[WIDTH-1:0] i3_mul1;
wire[WIDTH-1:0] i3_add1;
wire[WIDTH-1:0] i4_load;
wire[WIDTH-1:0] i5_add;
wire[WIDTH-1:0] i6_data_size1;
wire[WIDTH-1:0] i6_mul1;
wire[WIDTH-1:0] i6_add1;
wire[WIDTH-1:0] i7_load;
wire[WIDTH-1:0] i8_add;
wire[WIDTH-1:0] const3;
wire[WIDTH-1:0] i9_data_size1;
wire[WIDTH-1:0] i9_mul1;
wire[WIDTH-1:0] i9_add1;
wire[WIDTH-1:0] i10_load;
wire[WIDTH-1:0] const4;
wire[WIDTH-1:0] i11_add;
wire[WIDTH-1:0] i12_data_size1;
wire[WIDTH-1:0] i12_mul1;
wire[WIDTH-1:0] i12_add1;
wire[WIDTH-1:0] i13_load;
wire[WIDTH-1:0] i14_add;
wire[WIDTH-1:0] const5;
wire[WIDTH-1:0] i15_mul;
wire[WIDTH-1:0] i16_mul;
wire[WIDTH-1:0] i17_mul;
wire[WIDTH-1:0] i18_mul;
wire[WIDTH-1:0] i19_add;
wire[WIDTH-1:0] input0;
wire i20_icmp;
wire[WIDTH-1:0] const2_dup_1;
wire[WIDTH-1:0] const3_dup_1;
wire[WIDTH-1:0] const0_alu;
wire[WIDTH-1:0] const2_alu;
wire[WIDTH-1:0] i3_data_size1_alu;
wire[WIDTH-1:0] i3_mul1_alu;
wire[WIDTH-1:0] i3_add1_alu;
wire[WIDTH-1:0] i5_add_alu;
wire[WIDTH-1:0] i6_data_size1_alu;
wire[WIDTH-1:0] i6_mul1_alu;
wire[WIDTH-1:0] i6_add1_alu;
wire[WIDTH-1:0] i8_add_alu;
wire[WIDTH-1:0] const3_alu;
wire[WIDTH-1:0] i9_data_size1_alu;
wire[WIDTH-1:0] i9_mul1_alu;
wire[WIDTH-1:0] i9_add1_alu;
wire[WIDTH-1:0] const4_alu;
wire[WIDTH-1:0] i11_add_alu;
wire[WIDTH-1:0] i12_data_size1_alu;
wire[WIDTH-1:0] i12_mul1_alu;
wire[WIDTH-1:0] i12_add1_alu;
wire[WIDTH-1:0] i14_add_alu;
wire[WIDTH-1:0] const5_alu;
wire[WIDTH-1:0] i15_mul_alu;
wire[WIDTH-1:0] i16_mul_alu;
wire[WIDTH-1:0] i17_mul_alu;
wire[WIDTH-1:0] i18_mul_alu;
wire[WIDTH-1:0] i19_add_alu;
wire[WIDTH-1:0] i19_output_alu;
wire[WIDTH-1:0] const2_dup_1_alu;
wire[WIDTH-1:0] const3_dup_1_alu;
wire[WIDTH-1:0] i21_br;
wire[WIDTH-1:0] i19_output;


IO_WIDTH_1 inst_global_en(.from_fabric(), .in(), .to_fabric(global_en), .out());
IO_WIDTH_1 inst_global_rst(.from_fabric(), .in(), .to_fabric(global_rst), .out());

const_unit #(.ConfigBits(1)) inst_const0(.const_out(const0));
const_unit #(.ConfigBits(2560)) inst_const2(.const_out(const2));
const_unit #(.ConfigBits(4)) inst_i3_data_size1(.const_out(i3_data_size1));
ALU #(.ALU_func(mul_op)) inst_i3_mul1(.data_in1(i3_data_size1), .data_in2(i5_add), .data_in3(), .data_out(i3_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_mul1_reg(.reg_in(i3_mul1_alu), .reg_out(i3_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i3_add1(.data_in1(const2), .data_in2(i3_mul1), .data_in3(), .data_out(i3_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i3_add1_reg(.reg_in(i3_add1_alu), .reg_out(i3_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i4_load(.addr0(i3_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i4_load));
ALU #(.ALU_func(add_op)) inst_i5_add(.data_in1(const0), .data_in2(i5_add), .data_in3(), .data_out(i5_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i5_add_reg(.reg_in(i5_add_alu), .reg_out(i5_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i6_data_size1(.const_out(i6_data_size1));
ALU #(.ALU_func(mul_op)) inst_i6_mul1(.data_in1(i5_add), .data_in2(i6_data_size1), .data_in3(), .data_out(i6_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_mul1_reg(.reg_in(i6_mul1_alu), .reg_out(i6_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i6_add1(.data_in1(i6_mul1), .data_in2(const2_dup_1), .data_in3(), .data_out(i6_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i6_add1_reg(.reg_in(i6_add1_alu), .reg_out(i6_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i7_load(.addr0(i6_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i7_load));
ALU #(.ALU_func(add_op)) inst_i8_add(.data_in1(i4_load), .data_in2(i7_load), .data_in3(), .data_out(i8_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i8_add_reg(.reg_in(i8_add_alu), .reg_out(i8_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(2816)) inst_const3(.const_out(const3));
const_unit #(.ConfigBits(4)) inst_i9_data_size1(.const_out(i9_data_size1));
ALU #(.ALU_func(mul_op)) inst_i9_mul1(.data_in1(i9_data_size1), .data_in2(i5_add), .data_in3(), .data_out(i9_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_mul1_reg(.reg_in(i9_mul1_alu), .reg_out(i9_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i9_add1(.data_in1(const3), .data_in2(i9_mul1), .data_in3(), .data_out(i9_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i9_add1_reg(.reg_in(i9_add1_alu), .reg_out(i9_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i10_load(.addr0(i9_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i10_load));
const_unit #(.ConfigBits(3)) inst_const4(.const_out(const4));
ALU #(.ALU_func(add_op)) inst_i11_add(.data_in1(const4), .data_in2(i5_add), .data_in3(), .data_out(i11_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i11_add_reg(.reg_in(i11_add_alu), .reg_out(i11_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(4)) inst_i12_data_size1(.const_out(i12_data_size1));
ALU #(.ALU_func(mul_op)) inst_i12_mul1(.data_in1(i11_add), .data_in2(i12_data_size1), .data_in3(), .data_out(i12_mul1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_mul1_reg(.reg_in(i12_mul1_alu), .reg_out(i12_mul1), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i12_add1(.data_in1(i12_mul1), .data_in2(const3_dup_1), .data_in3(), .data_out(i12_add1_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i12_add1_reg(.reg_in(i12_add1_alu), .reg_out(i12_add1), .en(global_en), .rst(global_rst));
(* keep *)Mem #(.config_bits(0)) inst_i13_load(.addr0(i12_add1), .reset(global_rst), .write_data(), .write_en(), .read_data(i13_load));
ALU #(.ALU_func(add_op)) inst_i14_add(.data_in1(i10_load), .data_in2(i13_load), .data_in3(), .data_out(i14_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i14_add_reg(.reg_in(i14_add_alu), .reg_out(i14_add), .en(global_en), .rst(global_rst));
const_unit #(.ConfigBits(12)) inst_const5(.const_out(const5));
ALU #(.ALU_func(mul_op)) inst_i15_mul(.data_in1(i8_add), .data_in2(const5), .data_in3(), .data_out(i15_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i15_mul_reg(.reg_in(i15_mul_alu), .reg_out(i15_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i16_mul(.data_in1(i10_load), .data_in2(i15_mul), .data_in3(), .data_out(i16_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i16_mul_reg(.reg_in(i16_mul_alu), .reg_out(i16_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i17_mul(.data_in1(i13_load), .data_in2(i16_mul), .data_in3(), .data_out(i17_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i17_mul_reg(.reg_in(i17_mul_alu), .reg_out(i17_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(mul_op)) inst_i18_mul(.data_in1(i14_add), .data_in2(i17_mul), .data_in3(), .data_out(i18_mul_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i18_mul_reg(.reg_in(i18_mul_alu), .reg_out(i18_mul), .en(global_en), .rst(global_rst));
ALU #(.ALU_func(add_op)) inst_i19_add(.data_in1(i18_mul), .data_in2(i19_add), .data_in3(), .data_out(i19_add_alu));
reg_unit #(.tide_en(0), .tide_rst(0)) inst_i19_add_reg(.reg_in(i19_add_alu), .reg_out(i19_add), .en(global_en), .rst(global_rst));
(* keep *) IO inst_input0(.from_fabric(), .in(), .to_fabric(input0), .out());
compare #(.conf(0)) inst_i20_icmp(.A(i5_add), .B(input0), .Y(i20_icmp));
(* keep *) IO_WIDTH_1 inst_i21_br(.from_fabric(i20_icmp), .in(), .to_fabric(), .out());
(* keep *) IO inst_i19_output(.from_fabric(i19_add), .in(), .to_fabric(), .out());
const_unit #(.ConfigBits(2560)) inst_const2_dup_1(.const_out(const2_dup_1));
const_unit #(.ConfigBits(2816)) inst_const3_dup_1(.const_out(const3_dup_1));

endmodule
